magic
tech sky130A
magscale 1 2
timestamp 1669298116
<< metal1 >>
rect 71774 702992 71780 703044
rect 71832 703032 71838 703044
rect 72970 703032 72976 703044
rect 71832 703004 72976 703032
rect 71832 702992 71838 703004
rect 72970 702992 72976 703004
rect 73028 702992 73034 703044
rect 527266 700476 527272 700528
rect 527324 700516 527330 700528
rect 543458 700516 543464 700528
rect 527324 700488 543464 700516
rect 527324 700476 527330 700488
rect 543458 700476 543464 700488
rect 543516 700476 543522 700528
rect 495434 700408 495440 700460
rect 495492 700448 495498 700460
rect 510982 700448 510988 700460
rect 495492 700420 510988 700448
rect 495492 700408 495498 700420
rect 510982 700408 510988 700420
rect 511040 700408 511046 700460
rect 542354 700340 542360 700392
rect 542412 700380 542418 700392
rect 559650 700380 559656 700392
rect 542412 700352 559656 700380
rect 542412 700340 542418 700352
rect 559650 700340 559656 700352
rect 559708 700340 559714 700392
rect 342254 700272 342260 700324
rect 342312 700312 342318 700324
rect 348786 700312 348792 700324
rect 342312 700284 348792 700312
rect 342312 700272 342318 700284
rect 348786 700272 348792 700284
rect 348844 700272 348850 700324
rect 372614 700272 372620 700324
rect 372672 700312 372678 700324
rect 381170 700312 381176 700324
rect 372672 700284 381176 700312
rect 372672 700272 372678 700284
rect 381170 700272 381176 700284
rect 381228 700272 381234 700324
rect 387794 700272 387800 700324
rect 387852 700312 387858 700324
rect 397454 700312 397460 700324
rect 387852 700284 397460 700312
rect 387852 700272 387858 700284
rect 397454 700272 397460 700284
rect 397512 700272 397518 700324
rect 402974 700272 402980 700324
rect 403032 700312 403038 700324
rect 413646 700312 413652 700324
rect 403032 700284 413652 700312
rect 403032 700272 403038 700284
rect 413646 700272 413652 700284
rect 413704 700272 413710 700324
rect 419534 700272 419540 700324
rect 419592 700312 419598 700324
rect 429838 700312 429844 700324
rect 419592 700284 429844 700312
rect 419592 700272 419598 700284
rect 429838 700272 429844 700284
rect 429896 700272 429902 700324
rect 434714 700272 434720 700324
rect 434772 700312 434778 700324
rect 446122 700312 446128 700324
rect 434772 700284 446128 700312
rect 434772 700272 434778 700284
rect 446122 700272 446128 700284
rect 446180 700272 446186 700324
rect 449894 700272 449900 700324
rect 449952 700312 449958 700324
rect 462314 700312 462320 700324
rect 449952 700284 462320 700312
rect 449952 700272 449958 700284
rect 462314 700272 462320 700284
rect 462372 700272 462378 700324
rect 465074 700272 465080 700324
rect 465132 700312 465138 700324
rect 478506 700312 478512 700324
rect 465132 700284 478512 700312
rect 465132 700272 465138 700284
rect 478506 700272 478512 700284
rect 478564 700272 478570 700324
rect 480254 700272 480260 700324
rect 480312 700312 480318 700324
rect 494790 700312 494796 700324
rect 480312 700284 494796 700312
rect 480312 700272 480318 700284
rect 494790 700272 494796 700284
rect 494848 700272 494854 700324
rect 510614 700272 510620 700324
rect 510672 700312 510678 700324
rect 527174 700312 527180 700324
rect 510672 700284 527180 700312
rect 510672 700272 510678 700284
rect 527174 700272 527180 700284
rect 527232 700272 527238 700324
rect 557534 700272 557540 700324
rect 557592 700312 557598 700324
rect 575842 700312 575848 700324
rect 557592 700284 575848 700312
rect 557592 700272 557598 700284
rect 575842 700272 575848 700284
rect 575900 700272 575906 700324
rect 105446 699728 105452 699780
rect 105504 699768 105510 699780
rect 108298 699768 108304 699780
rect 105504 699740 108304 699768
rect 105504 699728 105510 699740
rect 108298 699728 108304 699740
rect 108356 699728 108362 699780
rect 121638 699660 121644 699712
rect 121696 699700 121702 699712
rect 124858 699700 124864 699712
rect 121696 699672 124864 699700
rect 121696 699660 121702 699672
rect 124858 699660 124864 699672
rect 124916 699660 124922 699712
rect 137830 699660 137836 699712
rect 137888 699700 137894 699712
rect 140038 699700 140044 699712
rect 137888 699672 140044 699700
rect 137888 699660 137894 699672
rect 140038 699660 140044 699672
rect 140096 699660 140102 699712
rect 154114 699660 154120 699712
rect 154172 699700 154178 699712
rect 156598 699700 156604 699712
rect 154172 699672 156604 699700
rect 154172 699660 154178 699672
rect 156598 699660 156604 699672
rect 156656 699660 156662 699712
rect 170306 699660 170312 699712
rect 170364 699700 170370 699712
rect 172514 699700 172520 699712
rect 170364 699672 172520 699700
rect 170364 699660 170370 699672
rect 172514 699660 172520 699672
rect 172572 699660 172578 699712
rect 186498 699660 186504 699712
rect 186556 699700 186562 699712
rect 189074 699700 189080 699712
rect 186556 699672 189080 699700
rect 186556 699660 186562 699672
rect 189074 699660 189080 699672
rect 189132 699660 189138 699712
rect 202782 699660 202788 699712
rect 202840 699700 202846 699712
rect 204254 699700 204260 699712
rect 202840 699672 204260 699700
rect 202840 699660 202846 699672
rect 204254 699660 204260 699672
rect 204312 699660 204318 699712
rect 249794 699660 249800 699712
rect 249852 699700 249858 699712
rect 251450 699700 251456 699712
rect 249852 699672 251456 699700
rect 249852 699660 249858 699672
rect 251450 699660 251456 699672
rect 251508 699660 251514 699712
rect 264974 699660 264980 699712
rect 265032 699700 265038 699712
rect 267642 699700 267648 699712
rect 265032 699672 267648 699700
rect 265032 699660 265038 699672
rect 267642 699660 267648 699672
rect 267700 699660 267706 699712
rect 280154 699660 280160 699712
rect 280212 699700 280218 699712
rect 283834 699700 283840 699712
rect 280212 699672 283840 699700
rect 280212 699660 280218 699672
rect 283834 699660 283840 699672
rect 283892 699660 283898 699712
rect 296714 699660 296720 699712
rect 296772 699700 296778 699712
rect 300118 699700 300124 699712
rect 296772 699672 300124 699700
rect 296772 699660 296778 699672
rect 300118 699660 300124 699672
rect 300176 699660 300182 699712
rect 311894 699660 311900 699712
rect 311952 699700 311958 699712
rect 316310 699700 316316 699712
rect 311952 699672 316316 699700
rect 311952 699660 311958 699672
rect 316310 699660 316316 699672
rect 316368 699660 316374 699712
rect 327074 699660 327080 699712
rect 327132 699700 327138 699712
rect 332502 699700 332508 699712
rect 327132 699672 332508 699700
rect 327132 699660 327138 699672
rect 332502 699660 332508 699672
rect 332560 699660 332566 699712
rect 569218 696940 569224 696992
rect 569276 696980 569282 696992
rect 580166 696980 580172 696992
rect 569276 696952 580172 696980
rect 569276 696940 569282 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 569310 683136 569316 683188
rect 569368 683176 569374 683188
rect 580166 683176 580172 683188
rect 569368 683148 580172 683176
rect 569368 683136 569374 683148
rect 580166 683136 580172 683148
rect 580224 683136 580230 683188
rect 6914 680960 6920 681012
rect 6972 681000 6978 681012
rect 19886 681000 19892 681012
rect 6972 680972 19892 681000
rect 6972 680960 6978 680972
rect 19886 680960 19892 680972
rect 19944 680960 19950 681012
rect 23474 680960 23480 681012
rect 23532 681000 23538 681012
rect 35250 681000 35256 681012
rect 23532 680972 35256 681000
rect 23532 680960 23538 680972
rect 35250 680960 35256 680972
rect 35308 680960 35314 681012
rect 40034 680960 40040 681012
rect 40092 681000 40098 681012
rect 50614 681000 50620 681012
rect 40092 680972 50620 681000
rect 40092 680960 40098 680972
rect 50614 680960 50620 680972
rect 50672 680960 50678 681012
rect 56594 680960 56600 681012
rect 56652 681000 56658 681012
rect 66254 681000 66260 681012
rect 56652 680972 66260 681000
rect 56652 680960 56658 680972
rect 66254 680960 66260 680972
rect 66312 680960 66318 681012
rect 71774 680960 71780 681012
rect 71832 681000 71838 681012
rect 81434 681000 81440 681012
rect 71832 680972 81440 681000
rect 71832 680960 71838 680972
rect 81434 680960 81440 680972
rect 81492 680960 81498 681012
rect 88334 680960 88340 681012
rect 88392 681000 88398 681012
rect 96706 681000 96712 681012
rect 88392 680972 96712 681000
rect 88392 680960 88398 680972
rect 96706 680960 96712 680972
rect 96764 680960 96770 681012
rect 140038 680756 140044 680808
rect 140096 680796 140102 680808
rect 142798 680796 142804 680808
rect 140096 680768 142804 680796
rect 140096 680756 140102 680768
rect 142798 680756 142804 680768
rect 142856 680756 142862 680808
rect 358538 680688 358544 680740
rect 358596 680728 358602 680740
rect 364334 680728 364340 680740
rect 358596 680700 364340 680728
rect 358596 680688 358602 680700
rect 364334 680688 364340 680700
rect 364392 680688 364398 680740
rect 108298 680552 108304 680604
rect 108356 680592 108362 680604
rect 112070 680592 112076 680604
rect 108356 680564 112076 680592
rect 108356 680552 108362 680564
rect 112070 680552 112076 680564
rect 112128 680552 112134 680604
rect 156598 680552 156604 680604
rect 156656 680592 156662 680604
rect 158162 680592 158168 680604
rect 156656 680564 158168 680592
rect 156656 680552 156662 680564
rect 158162 680552 158168 680564
rect 158220 680552 158226 680604
rect 218054 680552 218060 680604
rect 218112 680592 218118 680604
rect 219710 680592 219716 680604
rect 218112 680564 219716 680592
rect 218112 680552 218118 680564
rect 219710 680552 219716 680564
rect 219768 680552 219774 680604
rect 124858 680416 124864 680468
rect 124916 680456 124922 680468
rect 127434 680456 127440 680468
rect 124916 680428 127440 680456
rect 124916 680416 124922 680428
rect 127434 680416 127440 680428
rect 127492 680416 127498 680468
rect 569402 670692 569408 670744
rect 569460 670732 569466 670744
rect 580166 670732 580172 670744
rect 569460 670704 580172 670732
rect 569460 670692 569466 670704
rect 580166 670692 580172 670704
rect 580224 670692 580230 670744
rect 3418 670624 3424 670676
rect 3476 670664 3482 670676
rect 9398 670664 9404 670676
rect 3476 670636 9404 670664
rect 3476 670624 3482 670636
rect 9398 670624 9404 670636
rect 9456 670624 9462 670676
rect 3510 658180 3516 658232
rect 3568 658220 3574 658232
rect 9398 658220 9404 658232
rect 3568 658192 9404 658220
rect 3568 658180 3574 658192
rect 9398 658180 9404 658192
rect 9456 658180 9462 658232
rect 569218 656888 569224 656940
rect 569276 656928 569282 656940
rect 580166 656928 580172 656940
rect 569276 656900 580172 656928
rect 569276 656888 569282 656900
rect 580166 656888 580172 656900
rect 580224 656888 580230 656940
rect 3602 645804 3608 645856
rect 3660 645844 3666 645856
rect 9398 645844 9404 645856
rect 3660 645816 9404 645844
rect 3660 645804 3666 645816
rect 9398 645804 9404 645816
rect 9456 645804 9462 645856
rect 569310 643084 569316 643136
rect 569368 643124 569374 643136
rect 580166 643124 580172 643136
rect 569368 643096 580172 643124
rect 569368 643084 569374 643096
rect 580166 643084 580172 643096
rect 580224 643084 580230 643136
rect 3418 633360 3424 633412
rect 3476 633400 3482 633412
rect 8662 633400 8668 633412
rect 3476 633372 8668 633400
rect 3476 633360 3482 633372
rect 8662 633360 8668 633372
rect 8720 633360 8726 633412
rect 569218 630640 569224 630692
rect 569276 630680 569282 630692
rect 580166 630680 580172 630692
rect 569276 630652 580172 630680
rect 569276 630640 569282 630652
rect 580166 630640 580172 630652
rect 580224 630640 580230 630692
rect 3510 620916 3516 620968
rect 3568 620956 3574 620968
rect 8662 620956 8668 620968
rect 3568 620928 8668 620956
rect 3568 620916 3574 620928
rect 8662 620916 8668 620928
rect 8720 620916 8726 620968
rect 569310 616836 569316 616888
rect 569368 616876 569374 616888
rect 580166 616876 580172 616888
rect 569368 616848 580172 616876
rect 569368 616836 569374 616848
rect 580166 616836 580172 616848
rect 580224 616836 580230 616888
rect 3602 607928 3608 607980
rect 3660 607968 3666 607980
rect 9398 607968 9404 607980
rect 3660 607940 9404 607968
rect 3660 607928 3666 607940
rect 9398 607928 9404 607940
rect 9456 607928 9462 607980
rect 569402 603100 569408 603152
rect 569460 603140 569466 603152
rect 580166 603140 580172 603152
rect 569460 603112 580172 603140
rect 569460 603100 569466 603112
rect 580166 603100 580172 603112
rect 580224 603100 580230 603152
rect 3418 596096 3424 596148
rect 3476 596136 3482 596148
rect 9398 596136 9404 596148
rect 3476 596108 9404 596136
rect 3476 596096 3482 596108
rect 9398 596096 9404 596108
rect 9456 596096 9462 596148
rect 2774 592016 2780 592068
rect 2832 592056 2838 592068
rect 6270 592056 6276 592068
rect 2832 592028 6276 592056
rect 2832 592016 2838 592028
rect 6270 592016 6276 592028
rect 6328 592016 6334 592068
rect 569218 590656 569224 590708
rect 569276 590696 569282 590708
rect 579798 590696 579804 590708
rect 569276 590668 579804 590696
rect 569276 590656 569282 590668
rect 579798 590656 579804 590668
rect 579856 590656 579862 590708
rect 3510 585080 3516 585132
rect 3568 585120 3574 585132
rect 9398 585120 9404 585132
rect 3568 585092 9404 585120
rect 3568 585080 3574 585092
rect 9398 585080 9404 585092
rect 9456 585080 9462 585132
rect 2958 579640 2964 579692
rect 3016 579680 3022 579692
rect 6178 579680 6184 579692
rect 3016 579652 6184 579680
rect 3016 579640 3022 579652
rect 6178 579640 6184 579652
rect 6236 579640 6242 579692
rect 569310 576852 569316 576904
rect 569368 576892 569374 576904
rect 580166 576892 580172 576904
rect 569368 576864 580172 576892
rect 569368 576852 569374 576864
rect 580166 576852 580172 576864
rect 580224 576852 580230 576904
rect 6270 572636 6276 572688
rect 6328 572676 6334 572688
rect 8846 572676 8852 572688
rect 6328 572648 8852 572676
rect 6328 572636 6334 572648
rect 8846 572636 8852 572648
rect 8904 572636 8910 572688
rect 569218 563048 569224 563100
rect 569276 563088 569282 563100
rect 579798 563088 579804 563100
rect 569276 563060 579804 563088
rect 569276 563048 569282 563060
rect 579798 563048 579804 563060
rect 579856 563048 579862 563100
rect 6178 559784 6184 559836
rect 6236 559824 6242 559836
rect 9398 559824 9404 559836
rect 6236 559796 9404 559824
rect 6236 559784 6242 559796
rect 9398 559784 9404 559796
rect 9456 559784 9462 559836
rect 569310 550604 569316 550656
rect 569368 550644 569374 550656
rect 580166 550644 580172 550656
rect 569368 550616 580172 550644
rect 569368 550604 569374 550616
rect 580166 550604 580172 550616
rect 580224 550604 580230 550656
rect 3418 547816 3424 547868
rect 3476 547856 3482 547868
rect 9398 547856 9404 547868
rect 3476 547828 9404 547856
rect 3476 547816 3482 547828
rect 9398 547816 9404 547828
rect 9456 547816 9462 547868
rect 3418 539588 3424 539640
rect 3476 539628 3482 539640
rect 7650 539628 7656 539640
rect 3476 539600 7656 539628
rect 3476 539588 3482 539600
rect 7650 539588 7656 539600
rect 7708 539588 7714 539640
rect 569218 536800 569224 536852
rect 569276 536840 569282 536852
rect 580166 536840 580172 536852
rect 569276 536812 580172 536840
rect 569276 536800 569282 536812
rect 580166 536800 580172 536812
rect 580224 536800 580230 536852
rect 3510 535372 3516 535424
rect 3568 535412 3574 535424
rect 9398 535412 9404 535424
rect 3568 535384 9404 535412
rect 3568 535372 3574 535384
rect 9398 535372 9404 535384
rect 9456 535372 9462 535424
rect 3418 527144 3424 527196
rect 3476 527184 3482 527196
rect 7558 527184 7564 527196
rect 3476 527156 7564 527184
rect 3476 527144 3482 527156
rect 7558 527144 7564 527156
rect 7616 527144 7622 527196
rect 569310 524424 569316 524476
rect 569368 524464 569374 524476
rect 580166 524464 580172 524476
rect 569368 524436 580172 524464
rect 569368 524424 569374 524436
rect 580166 524424 580172 524436
rect 580224 524424 580230 524476
rect 3418 514768 3424 514820
rect 3476 514808 3482 514820
rect 8938 514808 8944 514820
rect 3476 514780 8944 514808
rect 3476 514768 3482 514780
rect 8938 514768 8944 514780
rect 8996 514768 9002 514820
rect 569218 510620 569224 510672
rect 569276 510660 569282 510672
rect 580166 510660 580172 510672
rect 569276 510632 580172 510660
rect 569276 510620 569282 510632
rect 580166 510620 580172 510632
rect 580224 510620 580230 510672
rect 3050 500964 3056 501016
rect 3108 501004 3114 501016
rect 9030 501004 9036 501016
rect 3108 500976 9036 501004
rect 3108 500964 3114 500976
rect 9030 500964 9036 500976
rect 9088 500964 9094 501016
rect 577498 496816 577504 496868
rect 577556 496856 577562 496868
rect 579890 496856 579896 496868
rect 577556 496828 579896 496856
rect 577556 496816 577562 496828
rect 579890 496816 579896 496828
rect 579948 496816 579954 496868
rect 3418 488656 3424 488708
rect 3476 488696 3482 488708
rect 8938 488696 8944 488708
rect 3476 488668 8944 488696
rect 3476 488656 3482 488668
rect 8938 488656 8944 488668
rect 8996 488656 9002 488708
rect 577590 484372 577596 484424
rect 577648 484412 577654 484424
rect 580626 484412 580632 484424
rect 577648 484384 580632 484412
rect 577648 484372 577654 484384
rect 580626 484372 580632 484384
rect 580684 484372 580690 484424
rect 569862 482944 569868 482996
rect 569920 482984 569926 482996
rect 577498 482984 577504 482996
rect 569920 482956 577504 482984
rect 569920 482944 569926 482956
rect 577498 482944 577504 482956
rect 577556 482944 577562 482996
rect 3418 475600 3424 475652
rect 3476 475640 3482 475652
rect 9030 475640 9036 475652
rect 3476 475612 9036 475640
rect 3476 475600 3482 475612
rect 9030 475600 9036 475612
rect 9088 475600 9094 475652
rect 576118 470568 576124 470620
rect 576176 470608 576182 470620
rect 579982 470608 579988 470620
rect 576176 470580 579988 470608
rect 576176 470568 576182 470580
rect 579982 470568 579988 470580
rect 580040 470568 580046 470620
rect 569862 470500 569868 470552
rect 569920 470540 569926 470552
rect 577590 470540 577596 470552
rect 569920 470512 577596 470540
rect 569920 470500 569926 470512
rect 577590 470500 577596 470512
rect 577648 470500 577654 470552
rect 3418 462544 3424 462596
rect 3476 462584 3482 462596
rect 8938 462584 8944 462596
rect 3476 462556 8944 462584
rect 3476 462544 3482 462556
rect 8938 462544 8944 462556
rect 8996 462544 9002 462596
rect 569862 457852 569868 457904
rect 569920 457892 569926 457904
rect 576118 457892 576124 457904
rect 569920 457864 576124 457892
rect 569920 457852 569926 457864
rect 576118 457852 576124 457864
rect 576176 457852 576182 457904
rect 2774 449420 2780 449472
rect 2832 449460 2838 449472
rect 6270 449460 6276 449472
rect 2832 449432 6276 449460
rect 2832 449420 2838 449432
rect 6270 449420 6276 449432
rect 6328 449420 6334 449472
rect 569126 445680 569132 445732
rect 569184 445720 569190 445732
rect 580258 445720 580264 445732
rect 569184 445692 580264 445720
rect 569184 445680 569190 445692
rect 580258 445680 580264 445692
rect 580316 445680 580322 445732
rect 6270 437384 6276 437436
rect 6328 437424 6334 437436
rect 9398 437424 9404 437436
rect 6328 437396 9404 437424
rect 6328 437384 6334 437396
rect 9398 437384 9404 437396
rect 9456 437384 9462 437436
rect 2958 436160 2964 436212
rect 3016 436200 3022 436212
rect 6178 436200 6184 436212
rect 3016 436172 6184 436200
rect 3016 436160 3022 436172
rect 6178 436160 6184 436172
rect 6236 436160 6242 436212
rect 569310 433236 569316 433288
rect 569368 433276 569374 433288
rect 580350 433276 580356 433288
rect 569368 433248 580356 433276
rect 569368 433236 569374 433248
rect 580350 433236 580356 433248
rect 580408 433236 580414 433288
rect 569218 430584 569224 430636
rect 569276 430624 569282 430636
rect 580166 430624 580172 430636
rect 569276 430596 580172 430624
rect 569276 430584 569282 430596
rect 580166 430584 580172 430596
rect 580224 430584 580230 430636
rect 6178 424396 6184 424448
rect 6236 424436 6242 424448
rect 9398 424436 9404 424448
rect 6236 424408 9404 424436
rect 6236 424396 6242 424408
rect 9398 424396 9404 424408
rect 9456 424396 9462 424448
rect 3418 423172 3424 423224
rect 3476 423212 3482 423224
rect 7558 423212 7564 423224
rect 3476 423184 7564 423212
rect 3476 423172 3482 423184
rect 7558 423172 7564 423184
rect 7616 423172 7622 423224
rect 569218 418140 569224 418192
rect 569276 418180 569282 418192
rect 580166 418180 580172 418192
rect 569276 418152 580172 418180
rect 569276 418140 569282 418152
rect 580166 418140 580172 418152
rect 580224 418140 580230 418192
rect 3142 409844 3148 409896
rect 3200 409884 3206 409896
rect 7558 409884 7564 409896
rect 3200 409856 7564 409884
rect 3200 409844 3206 409856
rect 7558 409844 7564 409856
rect 7616 409844 7622 409896
rect 574738 404336 574744 404388
rect 574796 404376 574802 404388
rect 580166 404376 580172 404388
rect 574796 404348 580172 404376
rect 574796 404336 574802 404348
rect 580166 404336 580172 404348
rect 580224 404336 580230 404388
rect 3418 397468 3424 397520
rect 3476 397508 3482 397520
rect 7558 397508 7564 397520
rect 3476 397480 7564 397508
rect 3476 397468 3482 397480
rect 7558 397468 7564 397480
rect 7616 397468 7622 397520
rect 569126 395768 569132 395820
rect 569184 395808 569190 395820
rect 574738 395808 574744 395820
rect 569184 395780 574744 395808
rect 569184 395768 569190 395780
rect 574738 395768 574744 395780
rect 574796 395768 574802 395820
rect 3418 383800 3424 383852
rect 3476 383840 3482 383852
rect 7558 383840 7564 383852
rect 3476 383812 7564 383840
rect 3476 383800 3482 383812
rect 7558 383800 7564 383812
rect 7616 383800 7622 383852
rect 569862 383596 569868 383648
rect 569920 383636 569926 383648
rect 578878 383636 578884 383648
rect 569920 383608 578884 383636
rect 569920 383596 569926 383608
rect 578878 383596 578884 383608
rect 578936 383596 578942 383648
rect 3418 371288 3424 371340
rect 3476 371328 3482 371340
rect 7558 371328 7564 371340
rect 3476 371300 7564 371328
rect 3476 371288 3482 371300
rect 7558 371288 7564 371300
rect 7616 371288 7622 371340
rect 569586 371152 569592 371204
rect 569644 371192 569650 371204
rect 578878 371192 578884 371204
rect 569644 371164 578884 371192
rect 569644 371152 569650 371164
rect 578878 371152 578884 371164
rect 578936 371152 578942 371204
rect 578234 364692 578240 364744
rect 578292 364732 578298 364744
rect 579614 364732 579620 364744
rect 578292 364704 579620 364732
rect 578292 364692 578298 364704
rect 579614 364692 579620 364704
rect 579672 364692 579678 364744
rect 569678 358708 569684 358760
rect 569736 358748 569742 358760
rect 578234 358748 578240 358760
rect 569736 358720 578240 358748
rect 569736 358708 569742 358720
rect 578234 358708 578240 358720
rect 578292 358708 578298 358760
rect 2774 357688 2780 357740
rect 2832 357728 2838 357740
rect 4798 357728 4804 357740
rect 2832 357700 4804 357728
rect 2832 357688 2838 357700
rect 4798 357688 4804 357700
rect 4856 357688 4862 357740
rect 4798 351840 4804 351892
rect 4856 351880 4862 351892
rect 8662 351880 8668 351892
rect 4856 351852 8668 351880
rect 4856 351840 4862 351852
rect 8662 351840 8668 351852
rect 8720 351840 8726 351892
rect 569678 346332 569684 346384
rect 569736 346372 569742 346384
rect 579522 346372 579528 346384
rect 569736 346344 579528 346372
rect 569736 346332 569742 346344
rect 579522 346332 579528 346344
rect 579580 346332 579586 346384
rect 4154 339396 4160 339448
rect 4212 339436 4218 339448
rect 9398 339436 9404 339448
rect 4212 339408 9404 339436
rect 4212 339396 4218 339408
rect 9398 339396 9404 339408
rect 9456 339396 9462 339448
rect 569218 338104 569224 338156
rect 569276 338144 569282 338156
rect 580166 338144 580172 338156
rect 569276 338116 580172 338144
rect 569276 338104 569282 338116
rect 580166 338104 580172 338116
rect 580224 338104 580230 338156
rect 3050 327020 3056 327072
rect 3108 327060 3114 327072
rect 9398 327060 9404 327072
rect 3108 327032 9404 327060
rect 3108 327020 3114 327032
rect 9398 327020 9404 327032
rect 9456 327020 9462 327072
rect 568666 321512 568672 321564
rect 568724 321552 568730 321564
rect 580166 321552 580172 321564
rect 568724 321524 580172 321552
rect 568724 321512 568730 321524
rect 580166 321512 580172 321524
rect 580224 321512 580230 321564
rect 3418 314576 3424 314628
rect 3476 314616 3482 314628
rect 9398 314616 9404 314628
rect 3476 314588 9404 314616
rect 3476 314576 3482 314588
rect 9398 314576 9404 314588
rect 9456 314576 9462 314628
rect 568942 311856 568948 311908
rect 569000 311896 569006 311908
rect 580166 311896 580172 311908
rect 569000 311868 580172 311896
rect 569000 311856 569006 311868
rect 580166 311856 580172 311868
rect 580224 311856 580230 311908
rect 3418 306144 3424 306196
rect 3476 306184 3482 306196
rect 9398 306184 9404 306196
rect 3476 306156 9404 306184
rect 3476 306144 3482 306156
rect 9398 306144 9404 306156
rect 9456 306144 9462 306196
rect 569862 295264 569868 295316
rect 569920 295304 569926 295316
rect 580350 295304 580356 295316
rect 569920 295276 580356 295304
rect 569920 295264 569926 295276
rect 580350 295264 580356 295276
rect 580408 295264 580414 295316
rect 3418 292544 3424 292596
rect 3476 292584 3482 292596
rect 9398 292584 9404 292596
rect 3476 292556 9404 292584
rect 3476 292544 3482 292556
rect 9398 292544 9404 292556
rect 9456 292544 9462 292596
rect 572714 284316 572720 284368
rect 572772 284356 572778 284368
rect 580166 284356 580172 284368
rect 572772 284328 580172 284356
rect 572772 284316 572778 284328
rect 580166 284316 580172 284328
rect 580224 284316 580230 284368
rect 569862 282684 569868 282736
rect 569920 282724 569926 282736
rect 572714 282724 572720 282736
rect 569920 282696 572720 282724
rect 569920 282684 569926 282696
rect 572714 282684 572720 282696
rect 572772 282684 572778 282736
rect 3418 279692 3424 279744
rect 3476 279732 3482 279744
rect 9214 279732 9220 279744
rect 3476 279704 9220 279732
rect 3476 279692 3482 279704
rect 9214 279692 9220 279704
rect 9272 279692 9278 279744
rect 572714 271872 572720 271924
rect 572772 271912 572778 271924
rect 579798 271912 579804 271924
rect 572772 271884 579804 271912
rect 572772 271872 572778 271884
rect 579798 271872 579804 271884
rect 579856 271872 579862 271924
rect 569310 270172 569316 270224
rect 569368 270212 569374 270224
rect 572714 270212 572720 270224
rect 569368 270184 572720 270212
rect 569368 270172 569374 270184
rect 572714 270172 572720 270184
rect 572772 270172 572778 270224
rect 3050 266364 3056 266416
rect 3108 266404 3114 266416
rect 9398 266404 9404 266416
rect 3108 266376 9404 266404
rect 3108 266364 3114 266376
rect 9398 266364 9404 266376
rect 9456 266364 9462 266416
rect 579706 258108 579712 258120
rect 579586 258080 579712 258108
rect 569126 258000 569132 258052
rect 569184 258040 569190 258052
rect 579586 258040 579614 258080
rect 579706 258068 579712 258080
rect 579764 258068 579770 258120
rect 569184 258012 579614 258040
rect 569184 258000 569190 258012
rect 3418 254056 3424 254108
rect 3476 254096 3482 254108
rect 9398 254096 9404 254108
rect 3476 254068 9404 254096
rect 3476 254056 3482 254068
rect 9398 254056 9404 254068
rect 9456 254056 9462 254108
rect 568666 244876 568672 244928
rect 568724 244916 568730 244928
rect 580166 244916 580172 244928
rect 568724 244888 580172 244916
rect 568724 244876 568730 244888
rect 580166 244876 580172 244888
rect 580224 244876 580230 244928
rect 3418 240864 3424 240916
rect 3476 240904 3482 240916
rect 9398 240904 9404 240916
rect 3476 240876 9404 240904
rect 3476 240864 3482 240876
rect 9398 240864 9404 240876
rect 9456 240864 9462 240916
rect 569862 232500 569868 232552
rect 569920 232540 569926 232552
rect 580166 232540 580172 232552
rect 569920 232512 580172 232540
rect 569920 232500 569926 232512
rect 580166 232500 580172 232512
rect 580224 232500 580230 232552
rect 3418 227944 3424 227996
rect 3476 227984 3482 227996
rect 8846 227984 8852 227996
rect 3476 227956 8852 227984
rect 3476 227944 3482 227956
rect 8846 227944 8852 227956
rect 8904 227944 8910 227996
rect 569494 219444 569500 219496
rect 569552 219484 569558 219496
rect 569552 219456 579614 219484
rect 569552 219444 569558 219456
rect 579586 219416 579614 219456
rect 580442 219416 580448 219428
rect 579586 219388 580448 219416
rect 580442 219376 580448 219388
rect 580500 219376 580506 219428
rect 3418 214956 3424 215008
rect 3476 214996 3482 215008
rect 8202 214996 8208 215008
rect 3476 214968 8208 214996
rect 3476 214956 3482 214968
rect 8202 214956 8208 214968
rect 8260 214956 8266 215008
rect 569862 207000 569868 207052
rect 569920 207040 569926 207052
rect 579522 207040 579528 207052
rect 569920 207012 579528 207040
rect 569920 207000 569926 207012
rect 579522 207000 579528 207012
rect 579580 207000 579586 207052
rect 3326 202172 3332 202224
rect 3384 202212 3390 202224
rect 8202 202212 8208 202224
rect 3384 202184 8208 202212
rect 3384 202172 3390 202184
rect 8202 202172 8208 202184
rect 8260 202172 8266 202224
rect 569310 194556 569316 194608
rect 569368 194596 569374 194608
rect 579522 194596 579528 194608
rect 569368 194568 579528 194596
rect 569368 194556 569374 194568
rect 579522 194556 579528 194568
rect 579580 194556 579586 194608
rect 3418 188844 3424 188896
rect 3476 188884 3482 188896
rect 8202 188884 8208 188896
rect 3476 188856 8208 188884
rect 3476 188844 3482 188856
rect 8202 188844 8208 188856
rect 8260 188844 8266 188896
rect 569402 182180 569408 182232
rect 569460 182220 569466 182232
rect 576854 182220 576860 182232
rect 569460 182192 576860 182220
rect 569460 182180 569466 182192
rect 576854 182180 576860 182192
rect 576912 182180 576918 182232
rect 576854 179324 576860 179376
rect 576912 179364 576918 179376
rect 580258 179364 580264 179376
rect 576912 179336 580264 179364
rect 576912 179324 576918 179336
rect 580258 179324 580264 179336
rect 580316 179324 580322 179376
rect 3418 176604 3424 176656
rect 3476 176644 3482 176656
rect 8202 176644 8208 176656
rect 3476 176616 8208 176644
rect 3476 176604 3482 176616
rect 8202 176604 8208 176616
rect 8260 176604 8266 176656
rect 569862 169736 569868 169788
rect 569920 169776 569926 169788
rect 577958 169776 577964 169788
rect 569920 169748 577964 169776
rect 569920 169736 569926 169748
rect 577958 169736 577964 169748
rect 578016 169736 578022 169788
rect 577958 166948 577964 167000
rect 578016 166988 578022 167000
rect 579982 166988 579988 167000
rect 578016 166960 579988 166988
rect 578016 166948 578022 166960
rect 579982 166948 579988 166960
rect 580040 166948 580046 167000
rect 3510 163344 3516 163396
rect 3568 163384 3574 163396
rect 8202 163384 8208 163396
rect 3568 163356 8208 163384
rect 3568 163344 3574 163356
rect 8202 163344 8208 163356
rect 8260 163344 8266 163396
rect 569862 157360 569868 157412
rect 569920 157400 569926 157412
rect 579522 157400 579528 157412
rect 569920 157372 579528 157400
rect 569920 157360 569926 157372
rect 579522 157360 579528 157372
rect 579580 157360 579586 157412
rect 3418 150356 3424 150408
rect 3476 150396 3482 150408
rect 8938 150396 8944 150408
rect 3476 150368 8944 150396
rect 3476 150356 3482 150368
rect 8938 150356 8944 150368
rect 8996 150356 9002 150408
rect 569862 144916 569868 144968
rect 569920 144956 569926 144968
rect 578878 144956 578884 144968
rect 569920 144928 578884 144956
rect 569920 144916 569926 144928
rect 578878 144916 578884 144928
rect 578936 144916 578942 144968
rect 3234 137912 3240 137964
rect 3292 137952 3298 137964
rect 8294 137952 8300 137964
rect 3292 137924 8300 137952
rect 3292 137912 3298 137924
rect 8294 137912 8300 137924
rect 8352 137912 8358 137964
rect 569862 132472 569868 132524
rect 569920 132512 569926 132524
rect 578234 132512 578240 132524
rect 569920 132484 578240 132512
rect 569920 132472 569926 132484
rect 578234 132472 578240 132484
rect 578292 132472 578298 132524
rect 4154 129752 4160 129804
rect 4212 129792 4218 129804
rect 9030 129792 9036 129804
rect 4212 129764 9036 129792
rect 4212 129752 4218 129764
rect 9030 129752 9036 129764
rect 9088 129752 9094 129804
rect 578234 126896 578240 126948
rect 578292 126936 578298 126948
rect 579614 126936 579620 126948
rect 578292 126908 579620 126936
rect 578292 126896 578298 126908
rect 579614 126896 579620 126908
rect 579672 126896 579678 126948
rect 4798 118668 4804 118720
rect 4856 118708 4862 118720
rect 9398 118708 9404 118720
rect 4856 118680 9404 118708
rect 4856 118668 4862 118680
rect 9398 118668 9404 118680
rect 9456 118668 9462 118720
rect 568666 118668 568672 118720
rect 568724 118708 568730 118720
rect 578878 118708 578884 118720
rect 568724 118680 578884 118708
rect 568724 118668 568730 118680
rect 578878 118668 578884 118680
rect 578936 118668 578942 118720
rect 2774 110712 2780 110764
rect 2832 110752 2838 110764
rect 4798 110752 4804 110764
rect 2832 110724 4804 110752
rect 2832 110712 2838 110724
rect 4798 110712 4804 110724
rect 4856 110712 4862 110764
rect 4798 106292 4804 106344
rect 4856 106332 4862 106344
rect 9398 106332 9404 106344
rect 4856 106304 9404 106332
rect 4856 106292 4862 106304
rect 9398 106292 9404 106304
rect 9456 106292 9462 106344
rect 569678 106292 569684 106344
rect 569736 106332 569742 106344
rect 578878 106332 578884 106344
rect 569736 106304 578884 106332
rect 569736 106292 569742 106304
rect 578878 106292 578884 106304
rect 578936 106292 578942 106344
rect 2774 97724 2780 97776
rect 2832 97764 2838 97776
rect 4798 97764 4804 97776
rect 2832 97736 4804 97764
rect 2832 97724 2838 97736
rect 4798 97724 4804 97736
rect 4856 97724 4862 97776
rect 569678 94392 569684 94444
rect 569736 94432 569742 94444
rect 576118 94432 576124 94444
rect 569736 94404 576124 94432
rect 569736 94392 569742 94404
rect 576118 94392 576124 94404
rect 576176 94392 576182 94444
rect 4798 93848 4804 93900
rect 4856 93888 4862 93900
rect 9398 93888 9404 93900
rect 4856 93860 9404 93888
rect 4856 93848 4862 93860
rect 9398 93848 9404 93860
rect 9456 93848 9462 93900
rect 576118 86912 576124 86964
rect 576176 86952 576182 86964
rect 580166 86952 580172 86964
rect 576176 86924 580172 86952
rect 576176 86912 576182 86924
rect 580166 86912 580172 86924
rect 580224 86912 580230 86964
rect 2774 85212 2780 85264
rect 2832 85252 2838 85264
rect 4798 85252 4804 85264
rect 2832 85224 4804 85252
rect 2832 85212 2838 85224
rect 4798 85212 4804 85224
rect 4856 85212 4862 85264
rect 569678 81404 569684 81456
rect 569736 81444 569742 81456
rect 578878 81444 578884 81456
rect 569736 81416 578884 81444
rect 569736 81404 569742 81416
rect 578878 81404 578884 81416
rect 578936 81404 578942 81456
rect 3418 71612 3424 71664
rect 3476 71652 3482 71664
rect 8938 71652 8944 71664
rect 3476 71624 8944 71652
rect 3476 71612 3482 71624
rect 8938 71612 8944 71624
rect 8996 71612 9002 71664
rect 569586 69028 569592 69080
rect 569644 69068 569650 69080
rect 578878 69068 578884 69080
rect 569644 69040 578884 69068
rect 569644 69028 569650 69040
rect 578878 69028 578884 69040
rect 578936 69028 578942 69080
rect 3142 59168 3148 59220
rect 3200 59208 3206 59220
rect 8938 59208 8944 59220
rect 3200 59180 8944 59208
rect 3200 59168 3206 59180
rect 8938 59168 8944 59180
rect 8996 59168 9002 59220
rect 4798 56584 4804 56636
rect 4856 56624 4862 56636
rect 8846 56624 8852 56636
rect 4856 56596 8852 56624
rect 4856 56584 4862 56596
rect 8846 56584 8852 56596
rect 8904 56584 8910 56636
rect 569126 56584 569132 56636
rect 569184 56624 569190 56636
rect 574738 56624 574744 56636
rect 569184 56596 574744 56624
rect 569184 56584 569190 56596
rect 574738 56584 574744 56596
rect 574796 56584 574802 56636
rect 574738 46860 574744 46912
rect 574796 46900 574802 46912
rect 580166 46900 580172 46912
rect 574796 46872 580172 46900
rect 574796 46860 574802 46872
rect 580166 46860 580172 46872
rect 580224 46860 580230 46912
rect 2774 45500 2780 45552
rect 2832 45540 2838 45552
rect 4798 45540 4804 45552
rect 2832 45512 4804 45540
rect 2832 45500 2838 45512
rect 4798 45500 4804 45512
rect 4856 45500 4862 45552
rect 4890 44140 4896 44192
rect 4948 44180 4954 44192
rect 9398 44180 9404 44192
rect 4948 44152 9404 44180
rect 4948 44140 4954 44152
rect 9398 44140 9404 44152
rect 9456 44140 9462 44192
rect 569862 44140 569868 44192
rect 569920 44180 569926 44192
rect 578878 44180 578884 44192
rect 569920 44152 578884 44180
rect 569920 44140 569926 44152
rect 578878 44140 578884 44152
rect 578936 44140 578942 44192
rect 2774 32852 2780 32904
rect 2832 32892 2838 32904
rect 4890 32892 4896 32904
rect 2832 32864 4896 32892
rect 2832 32852 2838 32864
rect 4890 32852 4896 32864
rect 4948 32852 4954 32904
rect 4798 31764 4804 31816
rect 4856 31804 4862 31816
rect 9030 31804 9036 31816
rect 4856 31776 9036 31804
rect 4856 31764 4862 31776
rect 9030 31764 9036 31776
rect 9088 31764 9094 31816
rect 569494 31764 569500 31816
rect 569552 31804 569558 31816
rect 578970 31804 578976 31816
rect 569552 31776 578976 31804
rect 569552 31764 569558 31776
rect 578970 31764 578976 31776
rect 579028 31764 579034 31816
rect 2774 20340 2780 20392
rect 2832 20380 2838 20392
rect 4798 20380 4804 20392
rect 2832 20352 4804 20380
rect 2832 20340 2838 20352
rect 4798 20340 4804 20352
rect 4856 20340 4862 20392
rect 569862 19320 569868 19372
rect 569920 19360 569926 19372
rect 578878 19360 578884 19372
rect 569920 19332 578884 19360
rect 569920 19320 569926 19332
rect 578878 19320 578884 19332
rect 578936 19320 578942 19372
rect 75914 9596 75920 9648
rect 75972 9636 75978 9648
rect 81710 9636 81716 9648
rect 75972 9608 81716 9636
rect 75972 9596 75978 9608
rect 81710 9596 81716 9608
rect 81768 9596 81774 9648
rect 122834 9596 122840 9648
rect 122892 9636 122898 9648
rect 123662 9636 123668 9648
rect 122892 9608 123668 9636
rect 122892 9596 122898 9608
rect 123662 9596 123668 9608
rect 123720 9596 123726 9648
rect 229094 9596 229100 9648
rect 229152 9636 229158 9648
rect 229646 9636 229652 9648
rect 229152 9608 229652 9636
rect 229152 9596 229158 9608
rect 229646 9596 229652 9608
rect 229704 9596 229710 9648
rect 448882 9596 448888 9648
rect 448940 9636 448946 9648
rect 462774 9636 462780 9648
rect 448940 9608 462780 9636
rect 448940 9596 448946 9608
rect 462774 9596 462780 9608
rect 462832 9596 462838 9648
rect 463234 9596 463240 9648
rect 463292 9636 463298 9648
rect 476298 9636 476304 9648
rect 463292 9608 476304 9636
rect 463292 9596 463298 9608
rect 476298 9596 476304 9608
rect 476356 9596 476362 9648
rect 478690 9596 478696 9648
rect 478748 9636 478754 9648
rect 491386 9636 491392 9648
rect 478748 9608 491392 9636
rect 478748 9596 478754 9608
rect 491386 9596 491392 9608
rect 491444 9596 491450 9648
rect 501874 9596 501880 9648
rect 501932 9636 501938 9648
rect 515950 9636 515956 9648
rect 501932 9608 515956 9636
rect 501932 9596 501938 9608
rect 515950 9596 515956 9608
rect 516008 9596 516014 9648
rect 518434 9596 518440 9648
rect 518492 9636 518498 9648
rect 532602 9636 532608 9648
rect 518492 9608 532608 9636
rect 518492 9596 518498 9608
rect 532602 9596 532608 9608
rect 532660 9596 532666 9648
rect 26326 9528 26332 9580
rect 26384 9568 26390 9580
rect 35342 9568 35348 9580
rect 26384 9540 35348 9568
rect 26384 9528 26390 9540
rect 35342 9528 35348 9540
rect 35400 9528 35406 9580
rect 35986 9528 35992 9580
rect 36044 9568 36050 9580
rect 44174 9568 44180 9580
rect 36044 9540 44180 9568
rect 36044 9528 36050 9540
rect 44174 9528 44180 9540
rect 44232 9528 44238 9580
rect 68646 9528 68652 9580
rect 68704 9568 68710 9580
rect 73982 9568 73988 9580
rect 68704 9540 73988 9568
rect 68704 9528 68710 9540
rect 73982 9528 73988 9540
rect 74040 9528 74046 9580
rect 78582 9528 78588 9580
rect 78640 9568 78646 9580
rect 82814 9568 82820 9580
rect 78640 9540 82820 9568
rect 78640 9528 78646 9540
rect 82814 9528 82820 9540
rect 82872 9528 82878 9580
rect 103606 9528 103612 9580
rect 103664 9568 103670 9580
rect 107102 9568 107108 9580
rect 103664 9540 107108 9568
rect 103664 9528 103670 9540
rect 107102 9528 107108 9540
rect 107160 9528 107166 9580
rect 109126 9528 109132 9580
rect 109184 9568 109190 9580
rect 112622 9568 112628 9580
rect 109184 9540 112628 9568
rect 109184 9528 109190 9540
rect 112622 9528 112628 9540
rect 112680 9528 112686 9580
rect 124214 9528 124220 9580
rect 124272 9568 124278 9580
rect 125870 9568 125876 9580
rect 124272 9540 125876 9568
rect 124272 9528 124278 9540
rect 125870 9528 125876 9540
rect 125928 9528 125934 9580
rect 203886 9528 203892 9580
rect 203944 9568 203950 9580
rect 206462 9568 206468 9580
rect 203944 9540 206468 9568
rect 203944 9528 203950 9540
rect 206462 9528 206468 9540
rect 206520 9528 206526 9580
rect 271138 9528 271144 9580
rect 271196 9568 271202 9580
rect 272426 9568 272432 9580
rect 271196 9540 272432 9568
rect 271196 9528 271202 9540
rect 272426 9528 272432 9540
rect 272484 9528 272490 9580
rect 321922 9528 321928 9580
rect 321980 9568 321986 9580
rect 324222 9568 324228 9580
rect 321980 9540 324228 9568
rect 321980 9528 321986 9540
rect 324222 9528 324228 9540
rect 324280 9528 324286 9580
rect 338482 9528 338488 9580
rect 338540 9568 338546 9580
rect 340782 9568 340788 9580
rect 338540 9540 340788 9568
rect 338540 9528 338546 9540
rect 340782 9528 340788 9540
rect 340840 9528 340846 9580
rect 381538 9528 381544 9580
rect 381596 9568 381602 9580
rect 382918 9568 382924 9580
rect 381596 9540 382924 9568
rect 381596 9528 381602 9540
rect 382918 9528 382924 9540
rect 382976 9528 382982 9580
rect 410242 9528 410248 9580
rect 410300 9568 410306 9580
rect 412358 9568 412364 9580
rect 410300 9540 412364 9568
rect 410300 9528 410306 9540
rect 412358 9528 412364 9540
rect 412416 9528 412422 9580
rect 445570 9528 445576 9580
rect 445628 9568 445634 9580
rect 459186 9568 459192 9580
rect 445628 9540 459192 9568
rect 445628 9528 445634 9540
rect 459186 9528 459192 9540
rect 459244 9528 459250 9580
rect 467650 9528 467656 9580
rect 467708 9568 467714 9580
rect 480622 9568 480628 9580
rect 467708 9540 480628 9568
rect 467708 9528 467714 9540
rect 480622 9528 480628 9540
rect 480680 9528 480686 9580
rect 482922 9528 482928 9580
rect 482980 9568 482986 9580
rect 496446 9568 496452 9580
rect 482980 9540 496452 9568
rect 482980 9528 482986 9540
rect 496446 9528 496452 9540
rect 496504 9528 496510 9580
rect 499482 9528 499488 9580
rect 499540 9568 499546 9580
rect 513190 9568 513196 9580
rect 499540 9540 513196 9568
rect 499540 9528 499546 9540
rect 513190 9528 513196 9540
rect 513248 9528 513254 9580
rect 516042 9528 516048 9580
rect 516100 9568 516106 9580
rect 528646 9568 528652 9580
rect 516100 9540 528652 9568
rect 516100 9528 516106 9540
rect 528646 9528 528652 9540
rect 528704 9528 528710 9580
rect 534994 9528 535000 9580
rect 535052 9568 535058 9580
rect 547874 9568 547880 9580
rect 535052 9540 547880 9568
rect 535052 9528 535058 9540
rect 547874 9528 547880 9540
rect 547932 9528 547938 9580
rect 17954 9460 17960 9512
rect 18012 9500 18018 9512
rect 24302 9500 24308 9512
rect 18012 9472 24308 9500
rect 18012 9460 18018 9472
rect 24302 9460 24308 9472
rect 24360 9460 24366 9512
rect 26418 9460 26424 9512
rect 26476 9500 26482 9512
rect 34514 9500 34520 9512
rect 26476 9472 34520 9500
rect 26476 9460 26482 9472
rect 34514 9460 34520 9472
rect 34572 9460 34578 9512
rect 34698 9460 34704 9512
rect 34756 9500 34762 9512
rect 41966 9500 41972 9512
rect 34756 9472 41972 9500
rect 34756 9460 34762 9472
rect 41966 9460 41972 9472
rect 42024 9460 42030 9512
rect 45738 9460 45744 9512
rect 45796 9500 45802 9512
rect 53006 9500 53012 9512
rect 45796 9472 53012 9500
rect 45796 9460 45802 9472
rect 53006 9460 53012 9472
rect 53064 9460 53070 9512
rect 68922 9460 68928 9512
rect 68980 9500 68986 9512
rect 73154 9500 73160 9512
rect 68980 9472 73160 9500
rect 68980 9460 68986 9472
rect 73154 9460 73160 9472
rect 73212 9460 73218 9512
rect 76098 9460 76104 9512
rect 76156 9500 76162 9512
rect 80606 9500 80612 9512
rect 76156 9472 80612 9500
rect 76156 9460 76162 9472
rect 80606 9460 80612 9472
rect 80664 9460 80670 9512
rect 84378 9460 84384 9512
rect 84436 9500 84442 9512
rect 88334 9500 88340 9512
rect 84436 9472 88340 9500
rect 84436 9460 84442 9472
rect 88334 9460 88340 9472
rect 88392 9460 88398 9512
rect 93854 9460 93860 9512
rect 93912 9500 93918 9512
rect 98270 9500 98276 9512
rect 93912 9472 98276 9500
rect 93912 9460 93918 9472
rect 98270 9460 98276 9472
rect 98328 9460 98334 9512
rect 98454 9460 98460 9512
rect 98512 9500 98518 9512
rect 101582 9500 101588 9512
rect 98512 9472 101588 9500
rect 98512 9460 98518 9472
rect 101582 9460 101588 9472
rect 101640 9460 101646 9512
rect 104986 9460 104992 9512
rect 105044 9500 105050 9512
rect 108206 9500 108212 9512
rect 105044 9472 108212 9500
rect 105044 9460 105050 9472
rect 108206 9460 108212 9472
rect 108264 9460 108270 9512
rect 109218 9460 109224 9512
rect 109276 9500 109282 9512
rect 111794 9500 111800 9512
rect 109276 9472 111800 9500
rect 109276 9460 109282 9472
rect 111794 9460 111800 9472
rect 111852 9460 111858 9512
rect 114554 9460 114560 9512
rect 114612 9500 114618 9512
rect 117314 9500 117320 9512
rect 114612 9472 117320 9500
rect 114612 9460 114618 9472
rect 117314 9460 117320 9472
rect 117372 9460 117378 9512
rect 118602 9460 118608 9512
rect 118660 9500 118666 9512
rect 119246 9500 119252 9512
rect 118660 9472 119252 9500
rect 118660 9460 118666 9472
rect 119246 9460 119252 9472
rect 119304 9460 119310 9512
rect 124122 9460 124128 9512
rect 124180 9500 124186 9512
rect 124766 9500 124772 9512
rect 124180 9472 124772 9500
rect 124180 9460 124186 9472
rect 124766 9460 124772 9472
rect 124824 9460 124830 9512
rect 129642 9460 129648 9512
rect 129700 9500 129706 9512
rect 130286 9500 130292 9512
rect 129700 9472 130292 9500
rect 129700 9460 129706 9472
rect 130286 9460 130292 9472
rect 130344 9460 130350 9512
rect 155954 9460 155960 9512
rect 156012 9500 156018 9512
rect 156782 9500 156788 9512
rect 156012 9472 156788 9500
rect 156012 9460 156018 9472
rect 156782 9460 156788 9472
rect 156840 9460 156846 9512
rect 161474 9460 161480 9512
rect 161532 9500 161538 9512
rect 162302 9500 162308 9512
rect 161532 9472 162308 9500
rect 161532 9460 161538 9472
rect 162302 9460 162308 9472
rect 162360 9460 162366 9512
rect 166994 9460 167000 9512
rect 167052 9500 167058 9512
rect 167822 9500 167828 9512
rect 167052 9472 167828 9500
rect 167052 9460 167058 9472
rect 167822 9460 167828 9472
rect 167880 9460 167886 9512
rect 172514 9460 172520 9512
rect 172572 9500 172578 9512
rect 173342 9500 173348 9512
rect 172572 9472 173348 9500
rect 172572 9460 172578 9472
rect 173342 9460 173348 9472
rect 173400 9460 173406 9512
rect 192018 9460 192024 9512
rect 192076 9500 192082 9512
rect 195422 9500 195428 9512
rect 192076 9472 195428 9500
rect 192076 9460 192082 9472
rect 195422 9460 195428 9472
rect 195480 9460 195486 9512
rect 200298 9460 200304 9512
rect 200356 9500 200362 9512
rect 203150 9500 203156 9512
rect 200356 9472 203156 9500
rect 200356 9460 200362 9472
rect 203150 9460 203156 9472
rect 203208 9460 203214 9512
rect 206186 9460 206192 9512
rect 206244 9500 206250 9512
rect 208670 9500 208676 9512
rect 206244 9472 208676 9500
rect 206244 9460 206250 9472
rect 208670 9460 208676 9472
rect 208728 9460 208734 9512
rect 209774 9460 209780 9512
rect 209832 9500 209838 9512
rect 211982 9500 211988 9512
rect 209832 9472 211988 9500
rect 209832 9460 209838 9472
rect 211982 9460 211988 9472
rect 212040 9460 212046 9512
rect 214466 9460 214472 9512
rect 214524 9500 214530 9512
rect 216674 9500 216680 9512
rect 214524 9472 216680 9500
rect 214524 9460 214530 9472
rect 216674 9460 216680 9472
rect 216732 9460 216738 9512
rect 216858 9460 216864 9512
rect 216916 9500 216922 9512
rect 218606 9500 218612 9512
rect 216916 9472 218612 9500
rect 216916 9460 216922 9472
rect 218606 9460 218612 9472
rect 218664 9460 218670 9512
rect 220446 9460 220452 9512
rect 220504 9500 220510 9512
rect 222194 9500 222200 9512
rect 220504 9472 222200 9500
rect 220504 9460 220510 9472
rect 222194 9460 222200 9472
rect 222252 9460 222258 9512
rect 222746 9460 222752 9512
rect 222804 9500 222810 9512
rect 224126 9500 224132 9512
rect 222804 9472 224132 9500
rect 222804 9460 222810 9472
rect 224126 9460 224132 9472
rect 224184 9460 224190 9512
rect 226334 9460 226340 9512
rect 226392 9500 226398 9512
rect 227714 9500 227720 9512
rect 226392 9472 227720 9500
rect 226392 9460 226398 9472
rect 227714 9460 227720 9472
rect 227772 9460 227778 9512
rect 235810 9460 235816 9512
rect 235868 9500 235874 9512
rect 236270 9500 236276 9512
rect 235868 9472 236276 9500
rect 235868 9460 235874 9472
rect 236270 9460 236276 9472
rect 236328 9460 236334 9512
rect 256602 9460 256608 9512
rect 256660 9500 256666 9512
rect 257062 9500 257068 9512
rect 256660 9472 257068 9500
rect 256660 9460 256666 9472
rect 257062 9460 257068 9472
rect 257120 9460 257126 9512
rect 258994 9460 259000 9512
rect 259052 9500 259058 9512
rect 259546 9500 259552 9512
rect 259052 9472 259552 9500
rect 259052 9460 259058 9472
rect 259546 9460 259552 9472
rect 259604 9460 259610 9512
rect 262122 9460 262128 9512
rect 262180 9500 262186 9512
rect 262950 9500 262956 9512
rect 262180 9472 262956 9500
rect 262180 9460 262186 9472
rect 262950 9460 262956 9472
rect 263008 9460 263014 9512
rect 264514 9460 264520 9512
rect 264572 9500 264578 9512
rect 265342 9500 265348 9512
rect 264572 9472 265348 9500
rect 264572 9460 264578 9472
rect 265342 9460 265348 9472
rect 265400 9460 265406 9512
rect 270034 9460 270040 9512
rect 270092 9500 270098 9512
rect 271230 9500 271236 9512
rect 270092 9472 271236 9500
rect 270092 9460 270098 9472
rect 271230 9460 271236 9472
rect 271288 9460 271294 9512
rect 273162 9460 273168 9512
rect 273220 9500 273226 9512
rect 274542 9500 274548 9512
rect 273220 9472 274548 9500
rect 273220 9460 273226 9472
rect 274542 9460 274548 9472
rect 274600 9460 274606 9512
rect 277762 9460 277768 9512
rect 277820 9500 277826 9512
rect 279510 9500 279516 9512
rect 277820 9472 279516 9500
rect 277820 9460 277826 9472
rect 279510 9460 279516 9472
rect 279568 9460 279574 9512
rect 279970 9460 279976 9512
rect 280028 9500 280034 9512
rect 281442 9500 281448 9512
rect 280028 9472 281448 9500
rect 280028 9460 280034 9472
rect 281442 9460 281448 9472
rect 281500 9460 281506 9512
rect 284202 9460 284208 9512
rect 284260 9500 284266 9512
rect 284662 9500 284668 9512
rect 284260 9472 284668 9500
rect 284260 9460 284266 9472
rect 284662 9460 284668 9472
rect 284720 9460 284726 9512
rect 287698 9460 287704 9512
rect 287756 9500 287762 9512
rect 288434 9500 288440 9512
rect 287756 9472 288440 9500
rect 287756 9460 287762 9472
rect 288434 9460 288440 9472
rect 288492 9460 288498 9512
rect 290918 9460 290924 9512
rect 290976 9500 290982 9512
rect 291654 9500 291660 9512
rect 290976 9472 291660 9500
rect 290976 9460 290982 9472
rect 291654 9460 291660 9472
rect 291712 9460 291718 9512
rect 293218 9460 293224 9512
rect 293276 9500 293282 9512
rect 294230 9500 294236 9512
rect 293276 9472 294236 9500
rect 293276 9460 293282 9472
rect 294230 9460 294236 9472
rect 294288 9460 294294 9512
rect 295242 9460 295248 9512
rect 295300 9500 295306 9512
rect 296254 9500 296260 9512
rect 295300 9472 296260 9500
rect 295300 9460 295306 9472
rect 296254 9460 296260 9472
rect 296312 9460 296318 9512
rect 297634 9460 297640 9512
rect 297692 9500 297698 9512
rect 298094 9500 298100 9512
rect 297692 9472 298100 9500
rect 297692 9460 297698 9472
rect 298094 9460 298100 9472
rect 298152 9460 298158 9512
rect 299842 9460 299848 9512
rect 299900 9500 299906 9512
rect 301314 9500 301320 9512
rect 299900 9472 301320 9500
rect 299900 9460 299906 9472
rect 301314 9460 301320 9472
rect 301372 9460 301378 9512
rect 303062 9460 303068 9512
rect 303120 9500 303126 9512
rect 304442 9500 304448 9512
rect 303120 9472 304448 9500
rect 303120 9460 303126 9472
rect 304442 9460 304448 9472
rect 304500 9460 304506 9512
rect 308674 9460 308680 9512
rect 308732 9500 308738 9512
rect 310422 9500 310428 9512
rect 308732 9472 310428 9500
rect 308732 9460 308738 9472
rect 310422 9460 310428 9472
rect 310480 9460 310486 9512
rect 311802 9460 311808 9512
rect 311860 9500 311866 9512
rect 313182 9500 313188 9512
rect 311860 9472 313188 9500
rect 311860 9460 311866 9472
rect 313182 9460 313188 9472
rect 313240 9460 313246 9512
rect 314194 9460 314200 9512
rect 314252 9500 314258 9512
rect 315850 9500 315856 9512
rect 314252 9472 315856 9500
rect 314252 9460 314258 9472
rect 315850 9460 315856 9472
rect 315908 9460 315914 9512
rect 319714 9460 319720 9512
rect 319772 9500 319778 9512
rect 321462 9500 321468 9512
rect 319772 9472 321468 9500
rect 319772 9460 319778 9472
rect 321462 9460 321468 9472
rect 321520 9460 321526 9512
rect 322842 9460 322848 9512
rect 322900 9500 322906 9512
rect 324130 9500 324136 9512
rect 322900 9472 324136 9500
rect 322900 9460 322906 9472
rect 324130 9460 324136 9472
rect 324188 9460 324194 9512
rect 325234 9460 325240 9512
rect 325292 9500 325298 9512
rect 326246 9500 326252 9512
rect 325292 9472 326252 9500
rect 325292 9460 325298 9472
rect 326246 9460 326252 9472
rect 326304 9460 326310 9512
rect 327442 9460 327448 9512
rect 327500 9500 327506 9512
rect 329742 9500 329748 9512
rect 327500 9472 329748 9500
rect 327500 9460 327506 9472
rect 329742 9460 329748 9472
rect 329800 9460 329806 9512
rect 330754 9460 330760 9512
rect 330812 9500 330818 9512
rect 332502 9500 332508 9512
rect 330812 9472 332508 9500
rect 330812 9460 330818 9472
rect 332502 9460 332508 9472
rect 332560 9460 332566 9512
rect 336274 9460 336280 9512
rect 336332 9500 336338 9512
rect 336734 9500 336740 9512
rect 336332 9472 336740 9500
rect 336332 9460 336338 9472
rect 336734 9460 336740 9472
rect 336792 9460 336798 9512
rect 339402 9460 339408 9512
rect 339460 9500 339466 9512
rect 340690 9500 340696 9512
rect 339460 9472 340696 9500
rect 339460 9460 339466 9472
rect 340690 9460 340696 9472
rect 340748 9460 340754 9512
rect 341794 9460 341800 9512
rect 341852 9500 341858 9512
rect 343542 9500 343548 9512
rect 341852 9472 343548 9500
rect 341852 9460 341858 9472
rect 343542 9460 343548 9472
rect 343600 9460 343606 9512
rect 347314 9460 347320 9512
rect 347372 9500 347378 9512
rect 349062 9500 349068 9512
rect 347372 9472 349068 9500
rect 347372 9460 347378 9472
rect 349062 9460 349068 9472
rect 349120 9460 349126 9512
rect 350442 9460 350448 9512
rect 350500 9500 350506 9512
rect 351086 9500 351092 9512
rect 350500 9472 351092 9500
rect 350500 9460 350506 9472
rect 351086 9460 351092 9472
rect 351144 9460 351150 9512
rect 351730 9460 351736 9512
rect 351788 9500 351794 9512
rect 353202 9500 353208 9512
rect 351788 9472 353208 9500
rect 351788 9460 351794 9472
rect 353202 9460 353208 9472
rect 353260 9460 353266 9512
rect 355042 9460 355048 9512
rect 355100 9500 355106 9512
rect 356146 9500 356152 9512
rect 355100 9472 356152 9500
rect 355100 9460 355106 9472
rect 356146 9460 356152 9472
rect 356204 9460 356210 9512
rect 357250 9460 357256 9512
rect 357308 9500 357314 9512
rect 358722 9500 358728 9512
rect 357308 9472 358728 9500
rect 357308 9460 357314 9472
rect 358722 9460 358728 9472
rect 358780 9460 358786 9512
rect 366082 9460 366088 9512
rect 366140 9500 366146 9512
rect 368382 9500 368388 9512
rect 366140 9472 368388 9500
rect 366140 9460 366146 9472
rect 368382 9460 368388 9472
rect 368440 9460 368446 9512
rect 370498 9460 370504 9512
rect 370556 9500 370562 9512
rect 372154 9500 372160 9512
rect 370556 9472 372160 9500
rect 370556 9460 370562 9472
rect 372154 9460 372160 9472
rect 372212 9460 372218 9512
rect 372522 9460 372528 9512
rect 372580 9500 372586 9512
rect 373350 9500 373356 9512
rect 372580 9472 373356 9500
rect 372580 9460 372586 9472
rect 373350 9460 373356 9472
rect 373408 9460 373414 9512
rect 376018 9460 376024 9512
rect 376076 9500 376082 9512
rect 378042 9500 378048 9512
rect 376076 9472 378048 9500
rect 376076 9460 376082 9472
rect 378042 9460 378048 9472
rect 378100 9460 378106 9512
rect 380434 9460 380440 9512
rect 380492 9500 380498 9512
rect 381722 9500 381728 9512
rect 380492 9472 381728 9500
rect 380492 9460 380498 9472
rect 381722 9460 381728 9472
rect 381780 9460 381786 9512
rect 385954 9460 385960 9512
rect 386012 9500 386018 9512
rect 387702 9500 387708 9512
rect 386012 9472 387708 9500
rect 386012 9460 386018 9472
rect 387702 9460 387708 9472
rect 387760 9460 387766 9512
rect 389082 9460 389088 9512
rect 389140 9500 389146 9512
rect 390462 9500 390468 9512
rect 389140 9472 390468 9500
rect 389140 9460 389146 9472
rect 390462 9460 390468 9472
rect 390520 9460 390526 9512
rect 391474 9460 391480 9512
rect 391532 9500 391538 9512
rect 392486 9500 392492 9512
rect 391532 9472 392492 9500
rect 391532 9460 391538 9472
rect 392486 9460 392492 9472
rect 392544 9460 392550 9512
rect 396994 9460 397000 9512
rect 397052 9500 397058 9512
rect 398742 9500 398748 9512
rect 397052 9472 398748 9500
rect 397052 9460 397058 9472
rect 398742 9460 398748 9472
rect 398800 9460 398806 9512
rect 400122 9460 400128 9512
rect 400180 9500 400186 9512
rect 401410 9500 401416 9512
rect 400180 9472 401416 9500
rect 400180 9460 400186 9472
rect 401410 9460 401416 9472
rect 401468 9460 401474 9512
rect 406930 9460 406936 9512
rect 406988 9500 406994 9512
rect 407390 9500 407396 9512
rect 406988 9472 407396 9500
rect 406988 9460 406994 9472
rect 407390 9460 407396 9472
rect 407448 9460 407454 9512
rect 408034 9460 408040 9512
rect 408092 9500 408098 9512
rect 408494 9500 408500 9512
rect 408092 9472 408500 9500
rect 408092 9460 408098 9472
rect 408494 9460 408500 9472
rect 408552 9460 408558 9512
rect 409138 9460 409144 9512
rect 409196 9500 409202 9512
rect 411162 9500 411168 9512
rect 409196 9472 411168 9500
rect 409196 9460 409202 9472
rect 411162 9460 411168 9472
rect 411220 9460 411226 9512
rect 413554 9460 413560 9512
rect 413612 9500 413618 9512
rect 414014 9500 414020 9512
rect 413612 9472 414020 9500
rect 413612 9460 413618 9472
rect 414014 9460 414020 9472
rect 414072 9460 414078 9512
rect 416498 9460 416504 9512
rect 416556 9500 416562 9512
rect 418062 9500 418068 9512
rect 416556 9472 418068 9500
rect 416556 9460 416562 9472
rect 418062 9460 418068 9472
rect 418120 9460 418126 9512
rect 419074 9460 419080 9512
rect 419132 9500 419138 9512
rect 420822 9500 420828 9512
rect 419132 9472 420828 9500
rect 419132 9460 419138 9472
rect 420822 9460 420828 9472
rect 420880 9460 420886 9512
rect 426802 9460 426808 9512
rect 426860 9500 426866 9512
rect 427814 9500 427820 9512
rect 426860 9472 427820 9500
rect 426860 9460 426866 9472
rect 427814 9460 427820 9472
rect 427872 9460 427878 9512
rect 444282 9460 444288 9512
rect 444340 9500 444346 9512
rect 458082 9500 458088 9512
rect 444340 9472 458088 9500
rect 444340 9460 444346 9472
rect 458082 9460 458088 9472
rect 458140 9460 458146 9512
rect 469858 9460 469864 9512
rect 469916 9500 469922 9512
rect 484302 9500 484308 9512
rect 469916 9472 484308 9500
rect 469916 9460 469922 9472
rect 484302 9460 484308 9472
rect 484360 9460 484366 9512
rect 486418 9460 486424 9512
rect 486476 9500 486482 9512
rect 499666 9500 499672 9512
rect 486476 9472 499672 9500
rect 486476 9460 486482 9472
rect 499666 9460 499672 9472
rect 499724 9460 499730 9512
rect 502978 9460 502984 9512
rect 503036 9500 503042 9512
rect 516502 9500 516508 9512
rect 503036 9472 516508 9500
rect 503036 9460 503042 9472
rect 516502 9460 516508 9472
rect 516560 9460 516566 9512
rect 528278 9460 528284 9512
rect 528336 9500 528342 9512
rect 540974 9500 540980 9512
rect 528336 9472 540980 9500
rect 528336 9460 528342 9472
rect 540974 9460 540980 9472
rect 541032 9460 541038 9512
rect 24946 9392 24952 9444
rect 25004 9432 25010 9444
rect 29822 9432 29828 9444
rect 25004 9404 29828 9432
rect 25004 9392 25010 9404
rect 29822 9392 29828 9404
rect 29880 9392 29886 9444
rect 33778 9392 33784 9444
rect 33836 9432 33842 9444
rect 40862 9432 40868 9444
rect 33836 9404 40868 9432
rect 33836 9392 33842 9404
rect 40862 9392 40868 9404
rect 40920 9392 40926 9444
rect 41322 9392 41328 9444
rect 41380 9432 41386 9444
rect 47486 9432 47492 9444
rect 41380 9404 47492 9432
rect 41380 9392 41386 9404
rect 47486 9392 47492 9404
rect 47544 9392 47550 9444
rect 52270 9392 52276 9444
rect 52328 9432 52334 9444
rect 58526 9432 58532 9444
rect 52328 9404 58532 9432
rect 52328 9392 52334 9404
rect 58526 9392 58532 9404
rect 58584 9392 58590 9444
rect 59262 9392 59268 9444
rect 59320 9432 59326 9444
rect 64046 9432 64052 9444
rect 59320 9404 64052 9432
rect 59320 9392 59326 9404
rect 64046 9392 64052 9404
rect 64104 9392 64110 9444
rect 66346 9392 66352 9444
rect 66404 9432 66410 9444
rect 71774 9432 71780 9444
rect 66404 9404 71780 9432
rect 66404 9392 66410 9404
rect 71774 9392 71780 9404
rect 71832 9392 71838 9444
rect 74626 9392 74632 9444
rect 74684 9432 74690 9444
rect 79502 9432 79508 9444
rect 74684 9404 79508 9432
rect 74684 9392 74690 9404
rect 79502 9392 79508 9404
rect 79560 9392 79566 9444
rect 89622 9392 89628 9444
rect 89680 9432 89686 9444
rect 92750 9432 92756 9444
rect 89680 9404 92756 9432
rect 89680 9392 89686 9404
rect 92750 9392 92756 9404
rect 92808 9392 92814 9444
rect 99466 9392 99472 9444
rect 99524 9432 99530 9444
rect 102686 9432 102692 9444
rect 99524 9404 102692 9432
rect 99524 9392 99530 9404
rect 102686 9392 102692 9404
rect 102744 9392 102750 9444
rect 106826 9392 106832 9444
rect 106884 9432 106890 9444
rect 109310 9432 109316 9444
rect 106884 9404 109316 9432
rect 106884 9392 106890 9404
rect 109310 9392 109316 9404
rect 109368 9392 109374 9444
rect 113266 9392 113272 9444
rect 113324 9432 113330 9444
rect 115934 9432 115940 9444
rect 113324 9404 115940 9432
rect 113324 9392 113330 9404
rect 115934 9392 115940 9404
rect 115992 9392 115998 9444
rect 117222 9392 117228 9444
rect 117280 9432 117286 9444
rect 118142 9432 118148 9444
rect 117280 9404 118148 9432
rect 117280 9392 117286 9404
rect 118142 9392 118148 9404
rect 118200 9392 118206 9444
rect 118694 9392 118700 9444
rect 118752 9432 118758 9444
rect 121454 9432 121460 9444
rect 118752 9404 121460 9432
rect 118752 9392 118758 9404
rect 121454 9392 121460 9404
rect 121512 9392 121518 9444
rect 128262 9392 128268 9444
rect 128320 9432 128326 9444
rect 129182 9432 129188 9444
rect 128320 9404 129188 9432
rect 128320 9392 128326 9404
rect 129182 9392 129188 9404
rect 129240 9392 129246 9444
rect 193214 9392 193220 9444
rect 193272 9432 193278 9444
rect 196526 9432 196532 9444
rect 193272 9404 196532 9432
rect 193272 9392 193278 9404
rect 196526 9392 196532 9404
rect 196584 9392 196590 9444
rect 205082 9392 205088 9444
rect 205140 9432 205146 9444
rect 207566 9432 207572 9444
rect 205140 9404 207572 9432
rect 205140 9392 205146 9404
rect 207566 9392 207572 9404
rect 207624 9392 207630 9444
rect 213362 9392 213368 9444
rect 213420 9432 213426 9444
rect 215294 9432 215300 9444
rect 213420 9404 215300 9432
rect 213420 9392 213426 9404
rect 215294 9392 215300 9404
rect 215352 9392 215358 9444
rect 215662 9392 215668 9444
rect 215720 9432 215726 9444
rect 217502 9432 217508 9444
rect 215720 9404 217508 9432
rect 215720 9392 215726 9404
rect 217502 9392 217508 9404
rect 217560 9392 217566 9444
rect 221550 9392 221556 9444
rect 221608 9432 221614 9444
rect 223022 9432 223028 9444
rect 221608 9404 223028 9432
rect 221608 9392 221614 9404
rect 223022 9392 223028 9404
rect 223080 9392 223086 9444
rect 225138 9392 225144 9444
rect 225196 9432 225202 9444
rect 226426 9432 226432 9444
rect 225196 9404 226432 9432
rect 225196 9392 225202 9404
rect 226426 9392 226432 9404
rect 226484 9392 226490 9444
rect 227530 9392 227536 9444
rect 227588 9432 227594 9444
rect 228542 9432 228548 9444
rect 227588 9404 228548 9432
rect 227588 9392 227594 9404
rect 228542 9392 228548 9404
rect 228600 9392 228606 9444
rect 272242 9392 272248 9444
rect 272300 9432 272306 9444
rect 273622 9432 273628 9444
rect 272300 9404 273628 9432
rect 272300 9392 272306 9404
rect 273622 9392 273628 9404
rect 273680 9392 273686 9444
rect 274450 9392 274456 9444
rect 274508 9432 274514 9444
rect 275922 9432 275928 9444
rect 274508 9404 275928 9432
rect 274508 9392 274514 9404
rect 275922 9392 275928 9404
rect 275980 9392 275986 9444
rect 281074 9392 281080 9444
rect 281132 9432 281138 9444
rect 282822 9432 282828 9444
rect 281132 9404 282828 9432
rect 281132 9392 281138 9404
rect 282822 9392 282828 9404
rect 282880 9392 282886 9444
rect 283282 9392 283288 9444
rect 283340 9432 283346 9444
rect 285398 9432 285404 9444
rect 283340 9404 285404 9432
rect 283340 9392 283346 9404
rect 285398 9392 285404 9404
rect 285456 9392 285462 9444
rect 289722 9392 289728 9444
rect 289780 9432 289786 9444
rect 291010 9432 291016 9444
rect 289780 9404 291016 9432
rect 289780 9392 289786 9404
rect 291010 9392 291016 9404
rect 291068 9392 291074 9444
rect 292114 9392 292120 9444
rect 292172 9432 292178 9444
rect 292942 9432 292948 9444
rect 292172 9404 292948 9432
rect 292172 9392 292178 9404
rect 292942 9392 292948 9404
rect 293000 9392 293006 9444
rect 294322 9392 294328 9444
rect 294380 9432 294386 9444
rect 295518 9432 295524 9444
rect 294380 9404 295524 9432
rect 294380 9392 294386 9404
rect 295518 9392 295524 9404
rect 295576 9392 295582 9444
rect 300762 9392 300768 9444
rect 300820 9432 300826 9444
rect 301866 9432 301872 9444
rect 300820 9404 301872 9432
rect 300820 9392 300826 9404
rect 301866 9392 301872 9404
rect 301924 9392 301930 9444
rect 302050 9392 302056 9444
rect 302108 9432 302114 9444
rect 303154 9432 303160 9444
rect 302108 9404 303160 9432
rect 302108 9392 302114 9404
rect 303154 9392 303160 9404
rect 303212 9392 303218 9444
rect 309778 9392 309784 9444
rect 309836 9432 309842 9444
rect 311526 9432 311532 9444
rect 309836 9404 311532 9432
rect 309836 9392 309842 9404
rect 311526 9392 311532 9404
rect 311584 9392 311590 9444
rect 324038 9392 324044 9444
rect 324096 9432 324102 9444
rect 325050 9432 325056 9444
rect 324096 9404 325056 9432
rect 324096 9392 324102 9404
rect 325050 9392 325056 9404
rect 325108 9392 325114 9444
rect 326338 9392 326344 9444
rect 326396 9432 326402 9444
rect 327074 9432 327080 9444
rect 326396 9404 327080 9432
rect 326396 9392 326402 9404
rect 327074 9392 327080 9404
rect 327132 9392 327138 9444
rect 328362 9392 328368 9444
rect 328420 9432 328426 9444
rect 329650 9432 329656 9444
rect 328420 9404 329656 9432
rect 328420 9392 328426 9404
rect 329650 9392 329656 9404
rect 329708 9392 329714 9444
rect 340598 9392 340604 9444
rect 340656 9432 340662 9444
rect 342162 9432 342168 9444
rect 340656 9404 342168 9432
rect 340656 9392 340662 9404
rect 342162 9392 342168 9404
rect 342220 9392 342226 9444
rect 349522 9392 349528 9444
rect 349580 9432 349586 9444
rect 351822 9432 351828 9444
rect 349580 9404 351828 9432
rect 349580 9392 349586 9404
rect 351822 9392 351828 9404
rect 351880 9392 351886 9444
rect 352834 9392 352840 9444
rect 352892 9432 352898 9444
rect 354490 9432 354496 9444
rect 352892 9404 354496 9432
rect 352892 9392 352898 9404
rect 354490 9392 354496 9404
rect 354548 9392 354554 9444
rect 358354 9392 358360 9444
rect 358412 9432 358418 9444
rect 360102 9432 360108 9444
rect 358412 9404 360108 9432
rect 358412 9392 358418 9404
rect 360102 9392 360108 9404
rect 360160 9392 360166 9444
rect 361482 9392 361488 9444
rect 361540 9432 361546 9444
rect 362862 9432 362868 9444
rect 361540 9404 362868 9432
rect 361540 9392 361546 9404
rect 362862 9392 362868 9404
rect 362920 9392 362926 9444
rect 367002 9392 367008 9444
rect 367060 9432 367066 9444
rect 368290 9432 368296 9444
rect 367060 9404 368296 9432
rect 367060 9392 367066 9404
rect 368290 9392 368296 9404
rect 368348 9392 368354 9444
rect 369394 9392 369400 9444
rect 369452 9432 369458 9444
rect 371142 9432 371148 9444
rect 369452 9404 371148 9432
rect 369452 9392 369458 9404
rect 371142 9392 371148 9404
rect 371200 9392 371206 9444
rect 374914 9392 374920 9444
rect 374972 9432 374978 9444
rect 375374 9432 375380 9444
rect 374972 9404 375380 9432
rect 374972 9392 374978 9404
rect 375374 9392 375380 9404
rect 375432 9392 375438 9444
rect 390370 9392 390376 9444
rect 390428 9432 390434 9444
rect 391842 9432 391848 9444
rect 390428 9404 391848 9432
rect 390428 9392 390434 9404
rect 391842 9392 391848 9404
rect 391900 9392 391906 9444
rect 401318 9392 401324 9444
rect 401376 9432 401382 9444
rect 402882 9432 402888 9444
rect 401376 9404 402888 9432
rect 401376 9392 401382 9404
rect 402882 9392 402888 9404
rect 402940 9392 402946 9444
rect 405642 9392 405648 9444
rect 405700 9432 405706 9444
rect 407022 9432 407028 9444
rect 405700 9404 407028 9432
rect 405700 9392 405706 9404
rect 407022 9392 407028 9404
rect 407080 9392 407086 9444
rect 410978 9392 410984 9444
rect 411036 9432 411042 9444
rect 412542 9432 412548 9444
rect 411036 9404 412548 9432
rect 411036 9392 411042 9404
rect 412542 9392 412548 9404
rect 412600 9392 412606 9444
rect 414658 9392 414664 9444
rect 414716 9432 414722 9444
rect 416682 9432 416688 9444
rect 414716 9404 416688 9432
rect 414716 9392 414722 9404
rect 416682 9392 416688 9404
rect 416740 9392 416746 9444
rect 417970 9392 417976 9444
rect 418028 9432 418034 9444
rect 419442 9432 419448 9444
rect 418028 9404 419448 9432
rect 418028 9392 418034 9404
rect 419442 9392 419448 9404
rect 419500 9392 419506 9444
rect 432322 9392 432328 9444
rect 432380 9432 432386 9444
rect 433334 9432 433340 9444
rect 432380 9404 433340 9432
rect 432380 9392 432386 9404
rect 433334 9392 433340 9404
rect 433392 9392 433398 9444
rect 437842 9392 437848 9444
rect 437900 9432 437906 9444
rect 438854 9432 438860 9444
rect 437900 9404 438860 9432
rect 437900 9392 437906 9404
rect 438854 9392 438860 9404
rect 438912 9392 438918 9444
rect 443362 9392 443368 9444
rect 443420 9432 443426 9444
rect 456886 9432 456892 9444
rect 443420 9404 456892 9432
rect 443420 9392 443426 9404
rect 456886 9392 456892 9404
rect 456944 9392 456950 9444
rect 457714 9392 457720 9444
rect 457772 9432 457778 9444
rect 471882 9432 471888 9444
rect 457772 9404 471888 9432
rect 457772 9392 457778 9404
rect 471882 9392 471888 9404
rect 471940 9392 471946 9444
rect 473170 9392 473176 9444
rect 473228 9432 473234 9444
rect 486326 9432 486332 9444
rect 473228 9404 486332 9432
rect 473228 9392 473234 9404
rect 486326 9392 486332 9404
rect 486384 9392 486390 9444
rect 489638 9392 489644 9444
rect 489696 9432 489702 9444
rect 503622 9432 503628 9444
rect 489696 9404 503628 9432
rect 489696 9392 489702 9404
rect 503622 9392 503628 9404
rect 503680 9392 503686 9444
rect 505002 9392 505008 9444
rect 505060 9432 505066 9444
rect 517606 9432 517612 9444
rect 505060 9404 517612 9432
rect 505060 9392 505066 9404
rect 517606 9392 517612 9404
rect 517664 9392 517670 9444
rect 522850 9392 522856 9444
rect 522908 9432 522914 9444
rect 536006 9432 536012 9444
rect 522908 9404 536012 9432
rect 522908 9392 522914 9404
rect 536006 9392 536012 9404
rect 536064 9392 536070 9444
rect 34882 9324 34888 9376
rect 34940 9364 34946 9376
rect 43070 9364 43076 9376
rect 34940 9336 43076 9364
rect 34940 9324 34946 9336
rect 43070 9324 43076 9336
rect 43128 9324 43134 9376
rect 43346 9324 43352 9376
rect 43404 9364 43410 9376
rect 49694 9364 49700 9376
rect 43404 9336 49700 9364
rect 43404 9324 43410 9336
rect 49694 9324 49700 9336
rect 49752 9324 49758 9376
rect 50982 9324 50988 9376
rect 51040 9364 51046 9376
rect 56594 9364 56600 9376
rect 51040 9336 56600 9364
rect 51040 9324 51046 9336
rect 56594 9324 56600 9336
rect 56652 9324 56658 9376
rect 64966 9324 64972 9376
rect 65024 9364 65030 9376
rect 70670 9364 70676 9376
rect 65024 9336 70676 9364
rect 65024 9324 65030 9336
rect 70670 9324 70676 9336
rect 70728 9324 70734 9376
rect 81526 9324 81532 9376
rect 81584 9364 81590 9376
rect 86126 9364 86132 9376
rect 81584 9336 86132 9364
rect 81584 9324 81590 9336
rect 86126 9324 86132 9336
rect 86184 9324 86190 9376
rect 95326 9324 95332 9376
rect 95384 9364 95390 9376
rect 99374 9364 99380 9376
rect 95384 9336 99380 9364
rect 95384 9324 95390 9336
rect 99374 9324 99380 9336
rect 99432 9324 99438 9376
rect 133874 9324 133880 9376
rect 133932 9364 133938 9376
rect 135806 9364 135812 9376
rect 133932 9336 135812 9364
rect 133932 9324 133938 9336
rect 135806 9324 135812 9336
rect 135864 9324 135870 9376
rect 143534 9324 143540 9376
rect 143592 9364 143598 9376
rect 144914 9364 144920 9376
rect 143592 9336 144920 9364
rect 143592 9324 143598 9336
rect 144914 9324 144920 9336
rect 144972 9324 144978 9376
rect 282178 9324 282184 9376
rect 282236 9364 282242 9376
rect 284202 9364 284208 9376
rect 282236 9336 284208 9364
rect 282236 9324 282242 9336
rect 284202 9324 284208 9336
rect 284260 9324 284266 9376
rect 316402 9324 316408 9376
rect 316460 9364 316466 9376
rect 317414 9364 317420 9376
rect 316460 9336 317420 9364
rect 316460 9324 316466 9336
rect 317414 9324 317420 9336
rect 317472 9324 317478 9376
rect 320818 9324 320824 9376
rect 320876 9364 320882 9376
rect 322842 9364 322848 9376
rect 320876 9336 322848 9364
rect 320876 9324 320882 9336
rect 322842 9324 322848 9336
rect 322900 9324 322906 9376
rect 331858 9324 331864 9376
rect 331916 9364 331922 9376
rect 333882 9364 333888 9376
rect 331916 9336 333888 9364
rect 331916 9324 331922 9336
rect 333882 9324 333888 9336
rect 333940 9324 333946 9376
rect 337378 9324 337384 9376
rect 337436 9364 337442 9376
rect 339402 9364 339408 9376
rect 337436 9336 339408 9364
rect 337436 9324 337442 9336
rect 339402 9324 339408 9336
rect 339460 9324 339466 9376
rect 377858 9324 377864 9376
rect 377916 9364 377922 9376
rect 379422 9364 379428 9376
rect 377916 9336 379428 9364
rect 377916 9324 377922 9336
rect 379422 9324 379428 9336
rect 379480 9324 379486 9376
rect 387058 9324 387064 9376
rect 387116 9364 387122 9376
rect 389082 9364 389088 9376
rect 387116 9336 389088 9364
rect 387116 9324 387122 9336
rect 389082 9324 389088 9336
rect 389140 9324 389146 9376
rect 393682 9324 393688 9376
rect 393740 9364 393746 9376
rect 394786 9364 394792 9376
rect 393740 9336 394792 9364
rect 393740 9324 393746 9336
rect 394786 9324 394792 9336
rect 394844 9324 394850 9376
rect 398098 9324 398104 9376
rect 398156 9364 398162 9376
rect 400122 9364 400128 9376
rect 398156 9336 400128 9364
rect 398156 9324 398162 9336
rect 400122 9324 400128 9336
rect 400180 9324 400186 9376
rect 433242 9324 433248 9376
rect 433300 9364 433306 9376
rect 446214 9364 446220 9376
rect 433300 9336 446220 9364
rect 433300 9324 433306 9336
rect 446214 9324 446220 9336
rect 446272 9324 446278 9376
rect 456518 9324 456524 9376
rect 456576 9364 456582 9376
rect 470502 9364 470508 9376
rect 456576 9336 470508 9364
rect 456576 9324 456582 9336
rect 470502 9324 470508 9336
rect 470560 9324 470566 9376
rect 476482 9324 476488 9376
rect 476540 9364 476546 9376
rect 490098 9364 490104 9376
rect 476540 9336 490104 9364
rect 476540 9324 476546 9336
rect 490098 9324 490104 9336
rect 490156 9324 490162 9376
rect 496354 9324 496360 9376
rect 496412 9364 496418 9376
rect 510154 9364 510160 9376
rect 496412 9336 510160 9364
rect 496412 9324 496418 9336
rect 510154 9324 510160 9336
rect 510212 9324 510218 9376
rect 514018 9324 514024 9376
rect 514076 9364 514082 9376
rect 527910 9364 527916 9376
rect 514076 9336 527916 9364
rect 514076 9324 514082 9336
rect 527910 9324 527916 9336
rect 527968 9324 527974 9376
rect 529474 9324 529480 9376
rect 529532 9364 529538 9376
rect 542354 9364 542360 9376
rect 529532 9336 542360 9364
rect 529532 9324 529538 9336
rect 542354 9324 542360 9336
rect 542412 9324 542418 9376
rect 23290 9256 23296 9308
rect 23348 9296 23354 9308
rect 28994 9296 29000 9308
rect 23348 9268 29000 9296
rect 23348 9256 23354 9268
rect 28994 9256 29000 9268
rect 29052 9256 29058 9308
rect 29914 9256 29920 9308
rect 29972 9296 29978 9308
rect 37550 9296 37556 9308
rect 29972 9268 37556 9296
rect 29972 9256 29978 9268
rect 37550 9256 37556 9268
rect 37608 9256 37614 9308
rect 46934 9256 46940 9308
rect 46992 9296 46998 9308
rect 54110 9296 54116 9308
rect 46992 9268 54116 9296
rect 46992 9256 46998 9268
rect 54110 9256 54116 9268
rect 54168 9256 54174 9308
rect 56686 9256 56692 9308
rect 56744 9296 56750 9308
rect 62942 9296 62948 9308
rect 56744 9268 62948 9296
rect 56744 9256 56750 9268
rect 62942 9256 62948 9268
rect 63000 9256 63006 9308
rect 63494 9256 63500 9308
rect 63552 9296 63558 9308
rect 69566 9296 69572 9308
rect 63552 9268 69572 9296
rect 63552 9256 63558 9268
rect 69566 9256 69572 9268
rect 69624 9256 69630 9308
rect 70946 9256 70952 9308
rect 71004 9296 71010 9308
rect 76190 9296 76196 9308
rect 71004 9268 76196 9296
rect 71004 9256 71010 9268
rect 76190 9256 76196 9268
rect 76248 9256 76254 9308
rect 79962 9256 79968 9308
rect 80020 9296 80026 9308
rect 84194 9296 84200 9308
rect 80020 9268 84200 9296
rect 80020 9256 80026 9268
rect 84194 9256 84200 9268
rect 84252 9256 84258 9308
rect 304258 9256 304264 9308
rect 304316 9296 304322 9308
rect 305730 9296 305736 9308
rect 304316 9268 305736 9296
rect 304316 9256 304322 9268
rect 305730 9256 305736 9268
rect 305788 9256 305794 9308
rect 342898 9256 342904 9308
rect 342956 9296 342962 9308
rect 343726 9296 343732 9308
rect 342956 9268 343732 9296
rect 342956 9256 342962 9268
rect 343726 9256 343732 9268
rect 343784 9256 343790 9308
rect 359458 9256 359464 9308
rect 359516 9296 359522 9308
rect 361482 9296 361488 9308
rect 359516 9268 361488 9296
rect 359516 9256 359522 9268
rect 361482 9256 361488 9268
rect 361540 9256 361546 9308
rect 403618 9256 403624 9308
rect 403676 9296 403682 9308
rect 404354 9296 404360 9308
rect 403676 9268 404360 9296
rect 403676 9256 403682 9268
rect 404354 9256 404360 9268
rect 404412 9256 404418 9308
rect 415762 9256 415768 9308
rect 415820 9296 415826 9308
rect 417970 9296 417976 9308
rect 415820 9268 417976 9296
rect 415820 9256 415826 9268
rect 417970 9256 417976 9268
rect 418028 9256 418034 9308
rect 429010 9256 429016 9308
rect 429068 9296 429074 9308
rect 429654 9296 429660 9308
rect 429068 9268 429660 9296
rect 429068 9256 429074 9268
rect 429654 9256 429660 9268
rect 429712 9256 429718 9308
rect 436738 9256 436744 9308
rect 436796 9296 436802 9308
rect 438670 9296 438676 9308
rect 436796 9268 438676 9296
rect 436796 9256 436802 9268
rect 438670 9256 438676 9268
rect 438728 9256 438734 9308
rect 438762 9256 438768 9308
rect 438820 9296 438826 9308
rect 452102 9296 452108 9308
rect 438820 9268 452108 9296
rect 438820 9256 438826 9268
rect 452102 9256 452108 9268
rect 452160 9256 452166 9308
rect 455322 9256 455328 9308
rect 455380 9296 455386 9308
rect 467834 9296 467840 9308
rect 455380 9268 467840 9296
rect 455380 9256 455386 9268
rect 467834 9256 467840 9268
rect 467892 9256 467898 9308
rect 482002 9256 482008 9308
rect 482060 9296 482066 9308
rect 495526 9296 495532 9308
rect 482060 9268 495532 9296
rect 482060 9256 482066 9268
rect 495526 9256 495532 9268
rect 495584 9256 495590 9308
rect 504082 9256 504088 9308
rect 504140 9296 504146 9308
rect 517514 9296 517520 9308
rect 504140 9268 517520 9296
rect 504140 9256 504146 9268
rect 517514 9256 517520 9268
rect 517572 9256 517578 9308
rect 519538 9256 519544 9308
rect 519596 9296 519602 9308
rect 533982 9296 533988 9308
rect 519596 9268 533988 9296
rect 519596 9256 519602 9268
rect 533982 9256 533988 9268
rect 534040 9256 534046 9308
rect 538122 9256 538128 9308
rect 538180 9296 538186 9308
rect 551830 9296 551836 9308
rect 538180 9268 551836 9296
rect 538180 9256 538186 9268
rect 551830 9256 551836 9268
rect 551888 9256 551894 9308
rect 25038 9188 25044 9240
rect 25096 9228 25102 9240
rect 33134 9228 33140 9240
rect 25096 9200 33140 9228
rect 25096 9188 25102 9200
rect 33134 9188 33140 9200
rect 33192 9188 33198 9240
rect 44358 9188 44364 9240
rect 44416 9228 44422 9240
rect 51902 9228 51908 9240
rect 44416 9200 51908 9228
rect 44416 9188 44422 9200
rect 51902 9188 51908 9200
rect 51960 9188 51966 9240
rect 53926 9188 53932 9240
rect 53984 9228 53990 9240
rect 60734 9228 60740 9240
rect 53984 9200 60740 9228
rect 53984 9188 53990 9200
rect 60734 9188 60740 9200
rect 60792 9188 60798 9240
rect 72418 9188 72424 9240
rect 72476 9228 72482 9240
rect 77294 9228 77300 9240
rect 72476 9200 77300 9228
rect 72476 9188 72482 9200
rect 77294 9188 77300 9200
rect 77352 9188 77358 9240
rect 92566 9188 92572 9240
rect 92624 9228 92630 9240
rect 96062 9228 96068 9240
rect 92624 9200 96068 9228
rect 92624 9188 92630 9200
rect 96062 9188 96068 9200
rect 96120 9188 96126 9240
rect 199102 9188 199108 9240
rect 199160 9228 199166 9240
rect 202046 9228 202052 9240
rect 199160 9200 202052 9228
rect 199160 9188 199166 9200
rect 202046 9188 202052 9200
rect 202104 9188 202110 9240
rect 275554 9188 275560 9240
rect 275612 9228 275618 9240
rect 277118 9228 277124 9240
rect 275612 9200 277124 9228
rect 275612 9188 275618 9200
rect 277118 9188 277124 9200
rect 277176 9188 277182 9240
rect 332962 9188 332968 9240
rect 333020 9228 333026 9240
rect 335078 9228 335084 9240
rect 333020 9200 335084 9228
rect 333020 9188 333026 9200
rect 335078 9188 335084 9200
rect 335136 9188 335142 9240
rect 344922 9188 344928 9240
rect 344980 9228 344986 9240
rect 345106 9228 345112 9240
rect 344980 9200 345112 9228
rect 344980 9188 344986 9200
rect 345106 9188 345112 9200
rect 345164 9188 345170 9240
rect 382642 9188 382648 9240
rect 382700 9228 382706 9240
rect 384390 9228 384396 9240
rect 382700 9200 384396 9228
rect 382700 9188 382706 9200
rect 384390 9188 384396 9200
rect 384448 9188 384454 9240
rect 442258 9188 442264 9240
rect 442316 9228 442322 9240
rect 455690 9228 455696 9240
rect 442316 9200 455696 9228
rect 442316 9188 442322 9200
rect 455690 9188 455696 9200
rect 455748 9188 455754 9240
rect 458818 9188 458824 9240
rect 458876 9228 458882 9240
rect 471974 9228 471980 9240
rect 458876 9200 471980 9228
rect 458876 9188 458882 9200
rect 471974 9188 471980 9200
rect 472032 9188 472038 9240
rect 475378 9188 475384 9240
rect 475436 9228 475442 9240
rect 488534 9228 488540 9240
rect 475436 9200 488540 9228
rect 475436 9188 475442 9200
rect 488534 9188 488540 9200
rect 488592 9188 488598 9240
rect 490834 9188 490840 9240
rect 490892 9228 490898 9240
rect 505002 9228 505008 9240
rect 490892 9200 505008 9228
rect 490892 9188 490898 9200
rect 505002 9188 505008 9200
rect 505060 9188 505066 9240
rect 507394 9188 507400 9240
rect 507452 9228 507458 9240
rect 520458 9228 520464 9240
rect 507452 9200 520464 9228
rect 507452 9188 507458 9200
rect 520458 9188 520464 9200
rect 520516 9188 520522 9240
rect 525058 9188 525064 9240
rect 525116 9228 525122 9240
rect 538858 9228 538864 9240
rect 525116 9200 538864 9228
rect 525116 9188 525122 9200
rect 538858 9188 538864 9200
rect 538916 9188 538922 9240
rect 17862 9120 17868 9172
rect 17920 9160 17926 9172
rect 18782 9160 18788 9172
rect 17920 9132 18788 9160
rect 17920 9120 17926 9132
rect 18782 9120 18788 9132
rect 18840 9120 18846 9172
rect 24026 9120 24032 9172
rect 24084 9160 24090 9172
rect 32030 9160 32036 9172
rect 24084 9132 32036 9160
rect 24084 9120 24090 9132
rect 32030 9120 32036 9132
rect 32088 9120 32094 9172
rect 32766 9120 32772 9172
rect 32824 9160 32830 9172
rect 40034 9160 40040 9172
rect 32824 9132 40040 9160
rect 32824 9120 32830 9132
rect 40034 9120 40040 9132
rect 40092 9120 40098 9172
rect 41506 9120 41512 9172
rect 41564 9160 41570 9172
rect 48590 9160 48596 9172
rect 41564 9132 48596 9160
rect 41564 9120 41570 9132
rect 48590 9120 48596 9132
rect 48648 9120 48654 9172
rect 49602 9120 49608 9172
rect 49660 9160 49666 9172
rect 55306 9160 55312 9172
rect 49660 9132 55312 9160
rect 49660 9120 49666 9132
rect 55306 9120 55312 9132
rect 55364 9120 55370 9172
rect 62666 9120 62672 9172
rect 62724 9160 62730 9172
rect 68462 9160 68468 9172
rect 62724 9132 68468 9160
rect 62724 9120 62730 9132
rect 68462 9120 68468 9132
rect 68520 9120 68526 9172
rect 87782 9120 87788 9172
rect 87840 9160 87846 9172
rect 91646 9160 91652 9172
rect 87840 9132 91652 9160
rect 87840 9120 87846 9132
rect 91646 9120 91652 9132
rect 91704 9120 91710 9172
rect 92474 9120 92480 9172
rect 92532 9160 92538 9172
rect 97166 9160 97172 9172
rect 92532 9132 97172 9160
rect 92532 9120 92538 9132
rect 97166 9120 97172 9132
rect 97224 9120 97230 9172
rect 111978 9120 111984 9172
rect 112036 9160 112042 9172
rect 114830 9160 114836 9172
rect 112036 9132 114836 9160
rect 112036 9120 112042 9132
rect 114830 9120 114836 9132
rect 114888 9120 114894 9172
rect 201494 9120 201500 9172
rect 201552 9160 201558 9172
rect 204254 9160 204260 9172
rect 201552 9132 204260 9160
rect 201552 9120 201558 9132
rect 204254 9120 204260 9132
rect 204312 9120 204318 9172
rect 210970 9120 210976 9172
rect 211028 9160 211034 9172
rect 213086 9160 213092 9172
rect 211028 9132 213092 9160
rect 211028 9120 211034 9132
rect 213086 9120 213092 9132
rect 213144 9120 213150 9172
rect 263410 9120 263416 9172
rect 263468 9160 263474 9172
rect 264146 9160 264152 9172
rect 263468 9132 264152 9160
rect 263468 9120 263474 9132
rect 264146 9120 264152 9132
rect 264204 9120 264210 9172
rect 268930 9120 268936 9172
rect 268988 9160 268994 9172
rect 270034 9160 270040 9172
rect 268988 9132 270040 9160
rect 268988 9120 268994 9132
rect 270034 9120 270040 9132
rect 270092 9120 270098 9172
rect 298738 9120 298744 9172
rect 298796 9160 298802 9172
rect 300670 9160 300676 9172
rect 298796 9132 300676 9160
rect 298796 9120 298802 9132
rect 300670 9120 300676 9132
rect 300728 9120 300734 9172
rect 318610 9120 318616 9172
rect 318668 9160 318674 9172
rect 320082 9160 320088 9172
rect 318668 9132 320088 9160
rect 318668 9120 318674 9132
rect 320082 9120 320088 9132
rect 320140 9120 320146 9172
rect 329558 9120 329564 9172
rect 329616 9160 329622 9172
rect 331122 9160 331128 9172
rect 329616 9132 331128 9160
rect 329616 9120 329622 9132
rect 331122 9120 331128 9132
rect 331180 9120 331186 9172
rect 425698 9120 425704 9172
rect 425756 9160 425762 9172
rect 427722 9160 427728 9172
rect 425756 9132 427728 9160
rect 425756 9120 425762 9132
rect 427722 9120 427728 9132
rect 427780 9120 427786 9172
rect 440050 9120 440056 9172
rect 440108 9160 440114 9172
rect 453298 9160 453304 9172
rect 440108 9132 453304 9160
rect 440108 9120 440114 9132
rect 453298 9120 453304 9132
rect 453356 9120 453362 9172
rect 462314 9160 462320 9172
rect 460906 9132 462320 9160
rect 23382 9052 23388 9104
rect 23440 9092 23446 9104
rect 30926 9092 30932 9104
rect 23440 9064 30932 9092
rect 23440 9052 23446 9064
rect 30926 9052 30932 9064
rect 30984 9052 30990 9104
rect 31662 9052 31668 9104
rect 31720 9092 31726 9104
rect 38654 9092 38660 9104
rect 31720 9064 38660 9092
rect 31720 9052 31726 9064
rect 38654 9052 38660 9064
rect 38712 9052 38718 9104
rect 82814 9052 82820 9104
rect 82872 9092 82878 9104
rect 87230 9092 87236 9104
rect 82872 9064 87236 9092
rect 82872 9052 82878 9064
rect 87230 9052 87236 9064
rect 87288 9052 87294 9104
rect 90174 9052 90180 9104
rect 90232 9092 90238 9104
rect 93946 9092 93952 9104
rect 90232 9064 93952 9092
rect 90232 9052 90238 9064
rect 93946 9052 93952 9064
rect 94004 9052 94010 9104
rect 373718 9052 373724 9104
rect 373776 9092 373782 9104
rect 374362 9092 374368 9104
rect 373776 9064 374368 9092
rect 373776 9052 373782 9064
rect 374362 9052 374368 9064
rect 374420 9052 374426 9104
rect 377122 9052 377128 9104
rect 377180 9092 377186 9104
rect 379238 9092 379244 9104
rect 377180 9064 379244 9092
rect 377180 9052 377186 9064
rect 379238 9052 379244 9064
rect 379296 9052 379302 9104
rect 427538 9052 427544 9104
rect 427596 9092 427602 9104
rect 440326 9092 440332 9104
rect 427596 9064 440332 9092
rect 427596 9052 427602 9064
rect 440326 9052 440332 9064
rect 440384 9052 440390 9104
rect 447778 9052 447784 9104
rect 447836 9092 447842 9104
rect 447836 9064 449756 9092
rect 447836 9052 447842 9064
rect 37274 8984 37280 9036
rect 37332 9024 37338 9036
rect 45554 9024 45560 9036
rect 37332 8996 45560 9024
rect 37332 8984 37338 8996
rect 45554 8984 45560 8996
rect 45612 8984 45618 9036
rect 73154 8984 73160 9036
rect 73212 9024 73218 9036
rect 78674 9024 78680 9036
rect 73212 8996 78680 9024
rect 73212 8984 73218 8996
rect 78674 8984 78680 8996
rect 78732 8984 78738 9036
rect 97166 8984 97172 9036
rect 97224 9024 97230 9036
rect 100754 9024 100760 9036
rect 97224 8996 100760 9024
rect 97224 8984 97230 8996
rect 100754 8984 100760 8996
rect 100812 8984 100818 9036
rect 102134 8984 102140 9036
rect 102192 9024 102198 9036
rect 106274 9024 106280 9036
rect 102192 8996 106280 9024
rect 102192 8984 102198 8996
rect 106274 8984 106280 8996
rect 106332 8984 106338 9036
rect 118050 8984 118056 9036
rect 118108 9024 118114 9036
rect 120350 9024 120356 9036
rect 118108 8996 120356 9024
rect 118108 8984 118114 8996
rect 120350 8984 120356 8996
rect 120408 8984 120414 9036
rect 212166 8984 212172 9036
rect 212224 9024 212230 9036
rect 214190 9024 214196 9036
rect 212224 8996 214196 9024
rect 212224 8984 212230 8996
rect 214190 8984 214196 8996
rect 214248 8984 214254 9036
rect 362770 8984 362776 9036
rect 362828 9024 362834 9036
rect 363322 9024 363328 9036
rect 362828 8996 363328 9024
rect 362828 8984 362834 8996
rect 363322 8984 363328 8996
rect 363380 8984 363386 9036
rect 364978 8984 364984 9036
rect 365036 9024 365042 9036
rect 365714 9024 365720 9036
rect 365036 8996 365720 9024
rect 365036 8984 365042 8996
rect 365714 8984 365720 8996
rect 365772 8984 365778 9036
rect 371602 8984 371608 9036
rect 371660 9024 371666 9036
rect 372614 9024 372620 9036
rect 371660 8996 372620 9024
rect 371660 8984 371666 8996
rect 372614 8984 372620 8996
rect 372672 8984 372678 9036
rect 435634 8984 435640 9036
rect 435692 9024 435698 9036
rect 448606 9024 448612 9036
rect 435692 8996 448612 9024
rect 435692 8984 435698 8996
rect 448606 8984 448612 8996
rect 448664 8984 448670 9036
rect 449728 9024 449756 9064
rect 449802 9052 449808 9104
rect 449860 9092 449866 9104
rect 460906 9092 460934 9132
rect 462314 9120 462320 9132
rect 462372 9120 462378 9172
rect 465442 9120 465448 9172
rect 465500 9160 465506 9172
rect 480162 9160 480168 9172
rect 465500 9132 480168 9160
rect 465500 9120 465506 9132
rect 480162 9120 480168 9132
rect 480220 9120 480226 9172
rect 480898 9120 480904 9172
rect 480956 9160 480962 9172
rect 495342 9160 495348 9172
rect 480956 9132 495348 9160
rect 480956 9120 480962 9132
rect 495342 9120 495348 9132
rect 495400 9120 495406 9172
rect 497458 9120 497464 9172
rect 497516 9160 497522 9172
rect 510706 9160 510712 9172
rect 497516 9132 510712 9160
rect 497516 9120 497522 9132
rect 510706 9120 510712 9132
rect 510764 9120 510770 9172
rect 517330 9120 517336 9172
rect 517388 9160 517394 9172
rect 530026 9160 530032 9172
rect 517388 9132 530032 9160
rect 517388 9120 517394 9132
rect 530026 9120 530032 9132
rect 530084 9120 530090 9172
rect 541618 9120 541624 9172
rect 541676 9160 541682 9172
rect 555418 9160 555424 9172
rect 541676 9132 555424 9160
rect 541676 9120 541682 9132
rect 555418 9120 555424 9132
rect 555476 9120 555482 9172
rect 449860 9064 460934 9092
rect 449860 9052 449866 9064
rect 464338 9052 464344 9104
rect 464396 9092 464402 9104
rect 478782 9092 478788 9104
rect 464396 9064 478788 9092
rect 464396 9052 464402 9064
rect 478782 9052 478788 9064
rect 478840 9052 478846 9104
rect 484210 9052 484216 9104
rect 484268 9092 484274 9104
rect 496906 9092 496912 9104
rect 484268 9064 496912 9092
rect 484268 9052 484274 9064
rect 496906 9052 496912 9064
rect 496964 9052 496970 9104
rect 500770 9052 500776 9104
rect 500828 9092 500834 9104
rect 514662 9092 514668 9104
rect 500828 9064 514668 9092
rect 500828 9052 500834 9064
rect 514662 9052 514668 9064
rect 514720 9052 514726 9104
rect 523954 9052 523960 9104
rect 524012 9092 524018 9104
rect 538030 9092 538036 9104
rect 524012 9064 538036 9092
rect 524012 9052 524018 9064
rect 538030 9052 538036 9064
rect 538088 9052 538094 9104
rect 544930 9052 544936 9104
rect 544988 9092 544994 9104
rect 557626 9092 557632 9104
rect 544988 9064 557632 9092
rect 544988 9052 544994 9064
rect 557626 9052 557632 9064
rect 557684 9052 557690 9104
rect 461578 9024 461584 9036
rect 449728 8996 461584 9024
rect 461578 8984 461584 8996
rect 461636 8984 461642 9036
rect 462130 8984 462136 9036
rect 462188 9024 462194 9036
rect 475102 9024 475108 9036
rect 462188 8996 475108 9024
rect 462188 8984 462194 8996
rect 475102 8984 475108 8996
rect 475160 8984 475166 9036
rect 477402 8984 477408 9036
rect 477460 9024 477466 9036
rect 490006 9024 490012 9036
rect 477460 8996 490012 9024
rect 477460 8984 477466 8996
rect 490006 8984 490012 8996
rect 490064 8984 490070 9036
rect 493042 8984 493048 9036
rect 493100 9024 493106 9036
rect 506474 9024 506480 9036
rect 493100 8996 506480 9024
rect 493100 8984 493106 8996
rect 506474 8984 506480 8996
rect 506532 8984 506538 9036
rect 520642 8984 520648 9036
rect 520700 9024 520706 9036
rect 534902 9024 534908 9036
rect 520700 8996 534908 9024
rect 520700 8984 520706 8996
rect 534902 8984 534908 8996
rect 534960 8984 534966 9036
rect 537202 8984 537208 9036
rect 537260 9024 537266 9036
rect 551922 9024 551928 9036
rect 537260 8996 551928 9024
rect 537260 8984 537266 8996
rect 551922 8984 551928 8996
rect 551980 8984 551986 9036
rect 15194 8916 15200 8968
rect 15252 8956 15258 8968
rect 20990 8956 20996 8968
rect 15252 8928 20996 8956
rect 15252 8916 15258 8928
rect 20990 8916 20996 8928
rect 21048 8916 21054 8968
rect 27614 8916 27620 8968
rect 27672 8956 27678 8968
rect 36446 8956 36452 8968
rect 27672 8928 36452 8956
rect 27672 8916 27678 8928
rect 36446 8916 36452 8928
rect 36504 8916 36510 8968
rect 43438 8916 43444 8968
rect 43496 8956 43502 8968
rect 51074 8956 51080 8968
rect 43496 8928 51080 8956
rect 43496 8916 43502 8928
rect 51074 8916 51080 8928
rect 51132 8916 51138 8968
rect 53098 8916 53104 8968
rect 53156 8956 53162 8968
rect 59630 8956 59636 8968
rect 53156 8928 59636 8956
rect 53156 8916 53162 8928
rect 59630 8916 59636 8928
rect 59688 8916 59694 8968
rect 60918 8916 60924 8968
rect 60976 8956 60982 8968
rect 67634 8956 67640 8968
rect 60976 8928 67640 8956
rect 60976 8916 60982 8928
rect 67634 8916 67640 8928
rect 67692 8916 67698 8968
rect 353938 8916 353944 8968
rect 353996 8956 354002 8968
rect 355042 8956 355048 8968
rect 353996 8928 355048 8956
rect 353996 8916 354002 8928
rect 355042 8916 355048 8928
rect 355100 8916 355106 8968
rect 402514 8916 402520 8968
rect 402572 8956 402578 8968
rect 403434 8956 403440 8968
rect 402572 8928 403440 8956
rect 402572 8916 402578 8928
rect 403434 8916 403440 8928
rect 403492 8916 403498 8968
rect 431218 8916 431224 8968
rect 431276 8956 431282 8968
rect 432230 8956 432236 8968
rect 431276 8928 432236 8956
rect 431276 8916 431282 8928
rect 432230 8916 432236 8928
rect 432288 8916 432294 8968
rect 434530 8916 434536 8968
rect 434588 8956 434594 8968
rect 447410 8956 447416 8968
rect 434588 8928 447416 8956
rect 434588 8916 434594 8928
rect 447410 8916 447416 8928
rect 447468 8916 447474 8968
rect 451090 8916 451096 8968
rect 451148 8956 451154 8968
rect 464982 8956 464988 8968
rect 451148 8928 464988 8956
rect 451148 8916 451154 8928
rect 464982 8916 464988 8928
rect 465040 8916 465046 8968
rect 470962 8916 470968 8968
rect 471020 8956 471026 8968
rect 484670 8956 484676 8968
rect 471020 8928 484676 8956
rect 471020 8916 471026 8928
rect 484670 8916 484676 8928
rect 484728 8916 484734 8968
rect 487522 8916 487528 8968
rect 487580 8956 487586 8968
rect 500954 8956 500960 8968
rect 487580 8928 500960 8956
rect 487580 8916 487586 8928
rect 500954 8916 500960 8928
rect 501012 8916 501018 8968
rect 510522 8916 510528 8968
rect 510580 8956 510586 8968
rect 524230 8956 524236 8968
rect 510580 8928 524236 8956
rect 510580 8916 510586 8928
rect 524230 8916 524236 8928
rect 524288 8916 524294 8968
rect 530578 8916 530584 8968
rect 530636 8956 530642 8968
rect 545022 8956 545028 8968
rect 530636 8928 545028 8956
rect 530636 8916 530642 8928
rect 545022 8916 545028 8928
rect 545080 8916 545086 8968
rect 547966 8916 547972 8968
rect 548024 8956 548030 8968
rect 568482 8956 568488 8968
rect 548024 8928 568488 8956
rect 548024 8916 548030 8928
rect 568482 8916 568488 8928
rect 568540 8916 568546 8968
rect 22094 8848 22100 8900
rect 22152 8888 22158 8900
rect 25406 8888 25412 8900
rect 22152 8860 25412 8888
rect 22152 8848 22158 8860
rect 25406 8848 25412 8860
rect 25464 8848 25470 8900
rect 55214 8848 55220 8900
rect 55272 8888 55278 8900
rect 62114 8888 62120 8900
rect 55272 8860 62120 8888
rect 55272 8848 55278 8860
rect 62114 8848 62120 8860
rect 62172 8848 62178 8900
rect 85574 8848 85580 8900
rect 85632 8888 85638 8900
rect 90542 8888 90548 8900
rect 85632 8860 90548 8888
rect 85632 8848 85638 8860
rect 90542 8848 90548 8860
rect 90600 8848 90606 8900
rect 126514 8848 126520 8900
rect 126572 8888 126578 8900
rect 128354 8888 128360 8900
rect 126572 8860 128360 8888
rect 126572 8848 126578 8860
rect 128354 8848 128360 8860
rect 128412 8848 128418 8900
rect 265618 8848 265624 8900
rect 265676 8888 265682 8900
rect 266538 8888 266544 8900
rect 265676 8860 266544 8888
rect 265676 8848 265682 8860
rect 266538 8848 266544 8860
rect 266596 8848 266602 8900
rect 285490 8848 285496 8900
rect 285548 8888 285554 8900
rect 286042 8888 286048 8900
rect 285548 8860 286048 8888
rect 285548 8848 285554 8860
rect 286042 8848 286048 8860
rect 286100 8848 286106 8900
rect 288802 8848 288808 8900
rect 288860 8888 288866 8900
rect 291102 8888 291108 8900
rect 288860 8860 291108 8888
rect 288860 8848 288866 8860
rect 291102 8848 291108 8860
rect 291160 8848 291166 8900
rect 313090 8848 313096 8900
rect 313148 8888 313154 8900
rect 314562 8888 314568 8900
rect 313148 8860 314568 8888
rect 313148 8848 313154 8860
rect 314562 8848 314568 8860
rect 314620 8848 314626 8900
rect 360562 8848 360568 8900
rect 360620 8888 360626 8900
rect 362770 8888 362776 8900
rect 360620 8860 362776 8888
rect 360620 8848 360626 8860
rect 362770 8848 362776 8860
rect 362828 8848 362834 8900
rect 388162 8848 388168 8900
rect 388220 8888 388226 8900
rect 390186 8888 390192 8900
rect 388220 8860 390192 8888
rect 388220 8848 388226 8860
rect 390186 8848 390192 8860
rect 390244 8848 390250 8900
rect 399202 8848 399208 8900
rect 399260 8888 399266 8900
rect 401502 8888 401508 8900
rect 399260 8860 401508 8888
rect 399260 8848 399266 8860
rect 401502 8848 401508 8860
rect 401560 8848 401566 8900
rect 471698 8848 471704 8900
rect 471756 8888 471762 8900
rect 485682 8888 485688 8900
rect 471756 8860 485688 8888
rect 471756 8848 471762 8860
rect 485682 8848 485688 8860
rect 485740 8848 485746 8900
rect 488442 8848 488448 8900
rect 488500 8888 488506 8900
rect 501046 8888 501052 8900
rect 488500 8860 501052 8888
rect 488500 8848 488506 8860
rect 501046 8848 501052 8860
rect 501104 8848 501110 8900
rect 506290 8848 506296 8900
rect 506348 8888 506354 8900
rect 518894 8888 518900 8900
rect 506348 8860 518900 8888
rect 506348 8848 506354 8860
rect 518894 8848 518900 8860
rect 518952 8848 518958 8900
rect 521562 8848 521568 8900
rect 521620 8888 521626 8900
rect 535362 8888 535368 8900
rect 521620 8860 535368 8888
rect 521620 8848 521626 8860
rect 535362 8848 535368 8860
rect 535420 8848 535426 8900
rect 363874 8780 363880 8832
rect 363932 8820 363938 8832
rect 364794 8820 364800 8832
rect 363932 8792 364800 8820
rect 363932 8780 363938 8792
rect 364794 8780 364800 8792
rect 364852 8780 364858 8832
rect 446674 8780 446680 8832
rect 446732 8820 446738 8832
rect 460382 8820 460388 8832
rect 446732 8792 460388 8820
rect 446732 8780 446738 8792
rect 460382 8780 460388 8792
rect 460440 8780 460446 8832
rect 460842 8780 460848 8832
rect 460900 8820 460906 8832
rect 474642 8820 474648 8832
rect 460900 8792 474648 8820
rect 460900 8780 460906 8792
rect 474642 8780 474648 8792
rect 474700 8780 474706 8832
rect 479794 8780 479800 8832
rect 479852 8820 479858 8832
rect 493962 8820 493968 8832
rect 479852 8792 493968 8820
rect 479852 8780 479858 8792
rect 493962 8780 493968 8792
rect 494020 8780 494026 8832
rect 508498 8780 508504 8832
rect 508556 8820 508562 8832
rect 522942 8820 522948 8832
rect 508556 8792 522948 8820
rect 508556 8780 508562 8792
rect 522942 8780 522948 8792
rect 523000 8780 523006 8832
rect 531498 8780 531504 8832
rect 531556 8820 531562 8832
rect 545758 8820 545764 8832
rect 531556 8792 545764 8820
rect 531556 8780 531562 8792
rect 545758 8780 545764 8792
rect 545816 8780 545822 8832
rect 108206 8712 108212 8764
rect 108264 8752 108270 8764
rect 110414 8752 110420 8764
rect 108264 8724 110420 8752
rect 108264 8712 108270 8724
rect 110414 8712 110420 8724
rect 110472 8712 110478 8764
rect 223942 8712 223948 8764
rect 224000 8752 224006 8764
rect 225230 8752 225236 8764
rect 224000 8724 225236 8752
rect 224000 8712 224006 8724
rect 225230 8712 225236 8724
rect 225288 8712 225294 8764
rect 231026 8712 231032 8764
rect 231084 8752 231090 8764
rect 231854 8752 231860 8764
rect 231084 8724 231860 8752
rect 231084 8712 231090 8724
rect 231854 8712 231860 8724
rect 231912 8712 231918 8764
rect 404722 8712 404728 8764
rect 404780 8752 404786 8764
rect 406102 8752 406108 8764
rect 404780 8724 406108 8752
rect 404780 8712 404786 8724
rect 406102 8712 406108 8724
rect 406160 8712 406166 8764
rect 420178 8712 420184 8764
rect 420236 8752 420242 8764
rect 420914 8752 420920 8764
rect 420236 8724 420920 8752
rect 420236 8712 420242 8724
rect 420914 8712 420920 8724
rect 420972 8712 420978 8764
rect 453206 8712 453212 8764
rect 453264 8752 453270 8764
rect 467466 8752 467472 8764
rect 453264 8724 467472 8752
rect 453264 8712 453270 8724
rect 467466 8712 467472 8724
rect 467524 8712 467530 8764
rect 474274 8712 474280 8764
rect 474332 8752 474338 8764
rect 487154 8752 487160 8764
rect 474332 8724 487160 8752
rect 474332 8712 474338 8724
rect 487154 8712 487160 8724
rect 487212 8712 487218 8764
rect 495250 8712 495256 8764
rect 495308 8752 495314 8764
rect 507854 8752 507860 8764
rect 495308 8724 507860 8752
rect 495308 8712 495314 8724
rect 507854 8712 507860 8724
rect 507912 8712 507918 8764
rect 511810 8712 511816 8764
rect 511868 8752 511874 8764
rect 525702 8752 525708 8764
rect 511868 8724 525708 8752
rect 511868 8712 511874 8724
rect 525702 8712 525708 8724
rect 525760 8712 525766 8764
rect 525794 8712 525800 8764
rect 525852 8752 525858 8764
rect 539686 8752 539692 8764
rect 525852 8724 539692 8752
rect 525852 8712 525858 8724
rect 539686 8712 539692 8724
rect 539744 8712 539750 8764
rect 344002 8644 344008 8696
rect 344060 8684 344066 8696
rect 345014 8684 345020 8696
rect 344060 8656 345020 8684
rect 344060 8644 344066 8656
rect 345014 8644 345020 8656
rect 345072 8644 345078 8696
rect 452194 8644 452200 8696
rect 452252 8684 452258 8696
rect 466270 8684 466276 8696
rect 452252 8656 466276 8684
rect 452252 8644 452258 8656
rect 466270 8644 466276 8656
rect 466328 8644 466334 8696
rect 468754 8644 468760 8696
rect 468812 8684 468818 8696
rect 481634 8684 481640 8696
rect 468812 8656 481640 8684
rect 468812 8644 468818 8656
rect 481634 8644 481640 8656
rect 481692 8644 481698 8696
rect 485314 8644 485320 8696
rect 485372 8684 485378 8696
rect 498194 8684 498200 8696
rect 485372 8656 498200 8684
rect 485372 8644 485378 8656
rect 498194 8644 498200 8656
rect 498252 8644 498258 8696
rect 512914 8644 512920 8696
rect 512972 8684 512978 8696
rect 526438 8684 526444 8696
rect 512972 8656 526444 8684
rect 512972 8644 512978 8656
rect 526438 8644 526444 8656
rect 526496 8644 526502 8696
rect 84286 8576 84292 8628
rect 84344 8616 84350 8628
rect 89714 8616 89720 8628
rect 84344 8588 89720 8616
rect 84344 8576 84350 8588
rect 89714 8576 89720 8588
rect 89772 8576 89778 8628
rect 348418 8576 348424 8628
rect 348476 8616 348482 8628
rect 350442 8616 350448 8628
rect 348476 8588 350448 8616
rect 348476 8576 348482 8588
rect 350442 8576 350448 8588
rect 350500 8576 350506 8628
rect 368198 8576 368204 8628
rect 368256 8616 368262 8628
rect 369762 8616 369768 8628
rect 368256 8588 369768 8616
rect 368256 8576 368262 8588
rect 369762 8576 369768 8588
rect 369820 8576 369826 8628
rect 424594 8576 424600 8628
rect 424652 8616 424658 8628
rect 426066 8616 426072 8628
rect 424652 8588 426072 8616
rect 424652 8576 424658 8588
rect 426066 8576 426072 8588
rect 426124 8576 426130 8628
rect 441154 8576 441160 8628
rect 441212 8616 441218 8628
rect 454494 8616 454500 8628
rect 441212 8588 454500 8616
rect 441212 8576 441218 8588
rect 454494 8576 454500 8588
rect 454552 8576 454558 8628
rect 466362 8576 466368 8628
rect 466420 8616 466426 8628
rect 478874 8616 478880 8628
rect 466420 8588 478880 8616
rect 466420 8576 466426 8588
rect 478874 8576 478880 8588
rect 478932 8576 478938 8628
rect 491938 8576 491944 8628
rect 491996 8616 492002 8628
rect 505554 8616 505560 8628
rect 491996 8588 505560 8616
rect 491996 8576 492002 8588
rect 505554 8576 505560 8588
rect 505612 8576 505618 8628
rect 515122 8576 515128 8628
rect 515180 8616 515186 8628
rect 528554 8616 528560 8628
rect 515180 8588 528560 8616
rect 515180 8576 515186 8588
rect 528554 8576 528560 8588
rect 528612 8576 528618 8628
rect 267642 8508 267648 8560
rect 267700 8548 267706 8560
rect 268838 8548 268844 8560
rect 267700 8520 268844 8548
rect 267700 8508 267706 8520
rect 268838 8508 268844 8520
rect 268896 8508 268902 8560
rect 306282 8508 306288 8560
rect 306340 8548 306346 8560
rect 306466 8548 306472 8560
rect 306340 8520 306472 8548
rect 306340 8508 306346 8520
rect 306466 8508 306472 8520
rect 306524 8508 306530 8560
rect 315298 8508 315304 8560
rect 315356 8548 315362 8560
rect 316034 8548 316040 8560
rect 315356 8520 316040 8548
rect 315356 8508 315362 8520
rect 316034 8508 316040 8520
rect 316092 8508 316098 8560
rect 383562 8508 383568 8560
rect 383620 8548 383626 8560
rect 383654 8548 383660 8560
rect 383620 8520 383660 8548
rect 383620 8508 383626 8520
rect 383654 8508 383660 8520
rect 383712 8508 383718 8560
rect 392578 8508 392584 8560
rect 392636 8548 392642 8560
rect 393314 8548 393320 8560
rect 392636 8520 393320 8548
rect 392636 8508 392642 8520
rect 393314 8508 393320 8520
rect 393372 8508 393378 8560
rect 421282 8508 421288 8560
rect 421340 8548 421346 8560
rect 423030 8548 423036 8560
rect 421340 8520 423036 8548
rect 421340 8508 421346 8520
rect 423030 8508 423036 8520
rect 423088 8508 423094 8560
rect 430114 8508 430120 8560
rect 430172 8548 430178 8560
rect 430942 8548 430948 8560
rect 430172 8520 430948 8548
rect 430172 8508 430178 8520
rect 430942 8508 430948 8520
rect 431000 8508 431006 8560
rect 454402 8508 454408 8560
rect 454460 8548 454466 8560
rect 468662 8548 468668 8560
rect 454460 8520 468668 8548
rect 454460 8508 454466 8520
rect 468662 8508 468668 8520
rect 468720 8508 468726 8560
rect 498562 8508 498568 8560
rect 498620 8548 498626 8560
rect 513282 8548 513288 8560
rect 498620 8520 513288 8548
rect 498620 8508 498626 8520
rect 513282 8508 513288 8520
rect 513340 8508 513346 8560
rect 207382 8440 207388 8492
rect 207440 8480 207446 8492
rect 209866 8480 209872 8492
rect 207440 8452 209872 8480
rect 207440 8440 207446 8452
rect 209866 8440 209872 8452
rect 209924 8440 209930 8492
rect 229830 8440 229836 8492
rect 229888 8480 229894 8492
rect 230750 8480 230756 8492
rect 229888 8452 230756 8480
rect 229888 8440 229894 8452
rect 230750 8440 230756 8452
rect 230808 8440 230814 8492
rect 310882 8440 310888 8492
rect 310940 8480 310946 8492
rect 312722 8480 312728 8492
rect 310940 8452 312728 8480
rect 310940 8440 310946 8452
rect 312722 8440 312728 8452
rect 312780 8440 312786 8492
rect 459922 8440 459928 8492
rect 459980 8480 459986 8492
rect 474550 8480 474556 8492
rect 459980 8452 474556 8480
rect 459980 8440 459986 8452
rect 474550 8440 474556 8452
rect 474608 8440 474614 8492
rect 493778 8440 493784 8492
rect 493836 8480 493842 8492
rect 506750 8480 506756 8492
rect 493836 8452 506756 8480
rect 493836 8440 493842 8452
rect 506750 8440 506756 8452
rect 506808 8440 506814 8492
rect 509602 8440 509608 8492
rect 509660 8480 509666 8492
rect 524322 8480 524328 8492
rect 509660 8452 524328 8480
rect 509660 8440 509666 8452
rect 524322 8440 524328 8452
rect 524380 8440 524386 8492
rect 60550 8372 60556 8424
rect 60608 8412 60614 8424
rect 65150 8412 65156 8424
rect 60608 8384 65156 8412
rect 60608 8372 60614 8384
rect 65150 8372 65156 8384
rect 65208 8372 65214 8424
rect 69934 8372 69940 8424
rect 69992 8412 69998 8424
rect 75086 8412 75092 8424
rect 69992 8384 75092 8412
rect 69992 8372 69998 8384
rect 75086 8372 75092 8384
rect 75144 8372 75150 8424
rect 100938 8372 100944 8424
rect 100996 8412 101002 8424
rect 103790 8412 103796 8424
rect 100996 8384 103796 8412
rect 100996 8372 101002 8384
rect 103790 8372 103796 8384
rect 103848 8372 103854 8424
rect 208578 8372 208584 8424
rect 208636 8412 208642 8424
rect 211154 8412 211160 8424
rect 208636 8384 211160 8412
rect 208636 8372 208642 8384
rect 211154 8372 211160 8384
rect 211212 8372 211218 8424
rect 219250 8372 219256 8424
rect 219308 8412 219314 8424
rect 220814 8412 220820 8424
rect 219308 8384 220820 8412
rect 219308 8372 219314 8384
rect 220814 8372 220820 8384
rect 220872 8372 220878 8424
rect 232222 8372 232228 8424
rect 232280 8412 232286 8424
rect 233234 8412 233240 8424
rect 232280 8384 233240 8412
rect 232280 8372 232286 8384
rect 233234 8372 233240 8384
rect 233292 8372 233298 8424
rect 257890 8372 257896 8424
rect 257948 8412 257954 8424
rect 258258 8412 258264 8424
rect 257948 8384 258264 8412
rect 257948 8372 257954 8384
rect 258258 8372 258264 8384
rect 258316 8372 258322 8424
rect 276658 8372 276664 8424
rect 276716 8412 276722 8424
rect 278314 8412 278320 8424
rect 276716 8384 278320 8412
rect 276716 8372 276722 8384
rect 278314 8372 278320 8384
rect 278372 8372 278378 8424
rect 379330 8372 379336 8424
rect 379388 8412 379394 8424
rect 380802 8412 380808 8424
rect 379388 8384 380808 8412
rect 379388 8372 379394 8384
rect 380802 8372 380808 8384
rect 380860 8372 380866 8424
rect 412450 8372 412456 8424
rect 412508 8412 412514 8424
rect 412634 8412 412640 8424
rect 412508 8384 412640 8412
rect 412508 8372 412514 8384
rect 412634 8372 412640 8384
rect 412692 8372 412698 8424
rect 13814 8304 13820 8356
rect 13872 8344 13878 8356
rect 16666 8344 16672 8356
rect 13872 8316 16672 8344
rect 13872 8304 13878 8316
rect 16666 8304 16672 8316
rect 16724 8304 16730 8356
rect 16758 8304 16764 8356
rect 16816 8344 16822 8356
rect 19886 8344 19892 8356
rect 16816 8316 19892 8344
rect 16816 8304 16822 8316
rect 19886 8304 19892 8316
rect 19944 8304 19950 8356
rect 39298 8304 39304 8356
rect 39356 8344 39362 8356
rect 46382 8344 46388 8356
rect 39356 8316 46388 8344
rect 39356 8304 39362 8316
rect 46382 8304 46388 8316
rect 46440 8304 46446 8356
rect 52086 8304 52092 8356
rect 52144 8344 52150 8356
rect 57422 8344 57428 8356
rect 52144 8316 57428 8344
rect 52144 8304 52150 8316
rect 57422 8304 57428 8316
rect 57480 8304 57486 8356
rect 59998 8304 60004 8356
rect 60056 8344 60062 8356
rect 66254 8344 66260 8356
rect 60056 8316 66260 8344
rect 60056 8304 60062 8316
rect 66254 8304 66260 8316
rect 66312 8304 66318 8356
rect 80514 8304 80520 8356
rect 80572 8344 80578 8356
rect 85022 8344 85028 8356
rect 80572 8316 85028 8344
rect 80572 8304 80578 8316
rect 85022 8304 85028 8316
rect 85080 8304 85086 8356
rect 91186 8304 91192 8356
rect 91244 8344 91250 8356
rect 95234 8344 95240 8356
rect 91244 8316 95240 8344
rect 91244 8304 91250 8316
rect 95234 8304 95240 8316
rect 95292 8304 95298 8356
rect 100846 8304 100852 8356
rect 100904 8344 100910 8356
rect 104894 8344 104900 8356
rect 100904 8316 104900 8344
rect 100904 8304 100910 8316
rect 104894 8304 104900 8316
rect 104952 8304 104958 8356
rect 110506 8304 110512 8356
rect 110564 8344 110570 8356
rect 113726 8344 113732 8356
rect 110564 8316 113732 8344
rect 110564 8304 110570 8316
rect 113726 8304 113732 8316
rect 113784 8304 113790 8356
rect 120166 8304 120172 8356
rect 120224 8344 120230 8356
rect 122926 8344 122932 8356
rect 120224 8316 122932 8344
rect 120224 8304 120230 8316
rect 122926 8304 122932 8316
rect 122984 8304 122990 8356
rect 197906 8304 197912 8356
rect 197964 8344 197970 8356
rect 200942 8344 200948 8356
rect 197964 8316 200948 8344
rect 197964 8304 197970 8316
rect 200942 8304 200948 8316
rect 201000 8304 201006 8356
rect 218054 8304 218060 8356
rect 218112 8344 218118 8356
rect 219710 8344 219716 8356
rect 218112 8316 219716 8344
rect 218112 8304 218118 8316
rect 219710 8304 219716 8316
rect 219768 8304 219774 8356
rect 238110 8304 238116 8356
rect 238168 8344 238174 8356
rect 238754 8344 238760 8356
rect 238168 8316 238760 8344
rect 238168 8304 238174 8316
rect 238754 8304 238760 8316
rect 238812 8304 238818 8356
rect 266722 8304 266728 8356
rect 266780 8344 266786 8356
rect 267734 8344 267740 8356
rect 266780 8316 267740 8344
rect 266780 8304 266786 8316
rect 267734 8304 267740 8316
rect 267792 8304 267798 8356
rect 286594 8304 286600 8356
rect 286652 8344 286658 8356
rect 287238 8344 287244 8356
rect 286652 8316 287244 8344
rect 286652 8304 286658 8316
rect 287238 8304 287244 8316
rect 287296 8304 287302 8356
rect 296530 8304 296536 8356
rect 296588 8344 296594 8356
rect 296714 8344 296720 8356
rect 296588 8316 296720 8344
rect 296588 8304 296594 8316
rect 296714 8304 296720 8316
rect 296772 8304 296778 8356
rect 305362 8304 305368 8356
rect 305420 8344 305426 8356
rect 306926 8344 306932 8356
rect 305420 8316 306932 8344
rect 305420 8304 305426 8316
rect 306926 8304 306932 8316
rect 306984 8304 306990 8356
rect 335170 8304 335176 8356
rect 335228 8344 335234 8356
rect 335354 8344 335360 8356
rect 335228 8316 335360 8344
rect 335228 8304 335234 8316
rect 335354 8304 335360 8316
rect 335412 8304 335418 8356
rect 422202 8304 422208 8356
rect 422260 8344 422266 8356
rect 422294 8344 422300 8356
rect 422260 8316 422300 8344
rect 422260 8304 422266 8316
rect 422294 8304 422300 8316
rect 422352 8304 422358 8356
rect 3418 6468 3424 6520
rect 3476 6508 3482 6520
rect 8938 6508 8944 6520
rect 3476 6480 8944 6508
rect 3476 6468 3482 6480
rect 8938 6468 8944 6480
rect 8996 6468 9002 6520
rect 5258 4088 5264 4140
rect 5316 4128 5322 4140
rect 15194 4128 15200 4140
rect 5316 4100 15200 4128
rect 5316 4088 5322 4100
rect 15194 4088 15200 4100
rect 15252 4088 15258 4140
rect 30098 4088 30104 4140
rect 30156 4128 30162 4140
rect 35986 4128 35992 4140
rect 30156 4100 35992 4128
rect 30156 4088 30162 4100
rect 35986 4088 35992 4100
rect 36044 4088 36050 4140
rect 39574 4088 39580 4140
rect 39632 4128 39638 4140
rect 45738 4128 45744 4140
rect 39632 4100 45744 4128
rect 39632 4088 39638 4100
rect 45738 4088 45744 4100
rect 45796 4088 45802 4140
rect 50154 4088 50160 4140
rect 50212 4128 50218 4140
rect 56686 4128 56692 4140
rect 50212 4100 56692 4128
rect 50212 4088 50218 4100
rect 56686 4088 56692 4100
rect 56744 4088 56750 4140
rect 58434 4088 58440 4140
rect 58492 4128 58498 4140
rect 64966 4128 64972 4140
rect 58492 4100 64972 4128
rect 58492 4088 58498 4100
rect 64966 4088 64972 4100
rect 65024 4088 65030 4140
rect 67910 4088 67916 4140
rect 67968 4128 67974 4140
rect 74626 4128 74632 4140
rect 67968 4100 74632 4128
rect 67968 4088 67974 4100
rect 74626 4088 74632 4100
rect 74684 4088 74690 4140
rect 79686 4088 79692 4140
rect 79744 4128 79750 4140
rect 85574 4128 85580 4140
rect 79744 4100 85580 4128
rect 79744 4088 79750 4100
rect 85574 4088 85580 4100
rect 85632 4088 85638 4140
rect 89162 4088 89168 4140
rect 89220 4128 89226 4140
rect 95234 4128 95240 4140
rect 89220 4100 95240 4128
rect 89220 4088 89226 4100
rect 95234 4088 95240 4100
rect 95292 4088 95298 4140
rect 97442 4088 97448 4140
rect 97500 4128 97506 4140
rect 103606 4128 103612 4140
rect 97500 4100 103612 4128
rect 97500 4088 97506 4100
rect 103606 4088 103612 4100
rect 103664 4088 103670 4140
rect 108114 4088 108120 4140
rect 108172 4128 108178 4140
rect 114554 4128 114560 4140
rect 108172 4100 114560 4128
rect 108172 4088 108178 4100
rect 114554 4088 114560 4100
rect 114612 4088 114618 4140
rect 116394 4088 116400 4140
rect 116452 4128 116458 4140
rect 124122 4128 124128 4140
rect 116452 4100 124128 4128
rect 116452 4088 116458 4100
rect 124122 4088 124128 4100
rect 124180 4088 124186 4140
rect 128170 4088 128176 4140
rect 128228 4128 128234 4140
rect 133874 4128 133880 4140
rect 128228 4100 133880 4128
rect 128228 4088 128234 4100
rect 133874 4088 133880 4100
rect 133932 4088 133938 4140
rect 137646 4088 137652 4140
rect 137704 4128 137710 4140
rect 143534 4128 143540 4140
rect 137704 4100 143540 4128
rect 137704 4088 137710 4100
rect 143534 4088 143540 4100
rect 143592 4088 143598 4140
rect 145926 4088 145932 4140
rect 145984 4128 145990 4140
rect 151814 4128 151820 4140
rect 145984 4100 151820 4128
rect 145984 4088 145990 4100
rect 151814 4088 151820 4100
rect 151872 4088 151878 4140
rect 157794 4088 157800 4140
rect 157852 4128 157858 4140
rect 162854 4128 162860 4140
rect 157852 4100 162860 4128
rect 157852 4088 157858 4100
rect 162854 4088 162860 4100
rect 162912 4088 162918 4140
rect 296254 4088 296260 4140
rect 296312 4128 296318 4140
rect 298462 4128 298468 4140
rect 296312 4100 298468 4128
rect 296312 4088 296318 4100
rect 298462 4088 298468 4100
rect 298520 4088 298526 4140
rect 324222 4088 324228 4140
rect 324280 4128 324286 4140
rect 326798 4128 326804 4140
rect 324280 4100 326804 4128
rect 324280 4088 324286 4100
rect 326798 4088 326804 4100
rect 326856 4088 326862 4140
rect 333882 4088 333888 4140
rect 333940 4128 333946 4140
rect 337470 4128 337476 4140
rect 333940 4100 337476 4128
rect 333940 4088 333946 4100
rect 337470 4088 337476 4100
rect 337528 4088 337534 4140
rect 342162 4088 342168 4140
rect 342220 4128 342226 4140
rect 346946 4128 346952 4140
rect 342220 4100 346952 4128
rect 342220 4088 342226 4100
rect 346946 4088 346952 4100
rect 347004 4088 347010 4140
rect 351822 4088 351828 4140
rect 351880 4128 351886 4140
rect 356330 4128 356336 4140
rect 351880 4100 356336 4128
rect 351880 4088 351886 4100
rect 356330 4088 356336 4100
rect 356388 4088 356394 4140
rect 358722 4088 358728 4140
rect 358780 4128 358786 4140
rect 364610 4128 364616 4140
rect 358780 4100 364616 4128
rect 358780 4088 358786 4100
rect 364610 4088 364616 4100
rect 364668 4088 364674 4140
rect 368290 4088 368296 4140
rect 368348 4128 368354 4140
rect 375282 4128 375288 4140
rect 368348 4100 375288 4128
rect 368348 4088 368354 4100
rect 375282 4088 375288 4100
rect 375340 4088 375346 4140
rect 387702 4088 387708 4140
rect 387760 4128 387766 4140
rect 395338 4128 395344 4140
rect 387760 4100 395344 4128
rect 387760 4088 387766 4100
rect 395338 4088 395344 4100
rect 395396 4088 395402 4140
rect 416682 4088 416688 4140
rect 416740 4128 416746 4140
rect 426158 4128 426164 4140
rect 416740 4100 426164 4128
rect 416740 4088 416746 4100
rect 426158 4088 426164 4100
rect 426216 4088 426222 4140
rect 506750 4088 506756 4140
rect 506808 4128 506814 4140
rect 511258 4128 511264 4140
rect 506808 4100 511264 4128
rect 506808 4088 506814 4100
rect 511258 4088 511264 4100
rect 511316 4088 511322 4140
rect 516502 4088 516508 4140
rect 516560 4128 516566 4140
rect 520734 4128 520740 4140
rect 516560 4100 520740 4128
rect 516560 4088 516566 4100
rect 520734 4088 520740 4100
rect 520792 4088 520798 4140
rect 525702 4088 525708 4140
rect 525760 4128 525766 4140
rect 530118 4128 530124 4140
rect 525760 4100 530124 4128
rect 525760 4088 525766 4100
rect 530118 4088 530124 4100
rect 530176 4088 530182 4140
rect 535362 4088 535368 4140
rect 535420 4128 535426 4140
rect 540790 4128 540796 4140
rect 535420 4100 540796 4128
rect 535420 4088 535426 4100
rect 540790 4088 540796 4100
rect 540848 4088 540854 4140
rect 542722 4088 542728 4140
rect 542780 4128 542786 4140
rect 563238 4128 563244 4140
rect 542780 4100 563244 4128
rect 542780 4088 542786 4100
rect 563238 4088 563244 4100
rect 563296 4088 563302 4140
rect 14734 4020 14740 4072
rect 14792 4060 14798 4072
rect 24946 4060 24952 4072
rect 14792 4032 24952 4060
rect 14792 4020 14798 4032
rect 24946 4020 24952 4032
rect 25004 4020 25010 4072
rect 53742 4020 53748 4072
rect 53800 4060 53806 4072
rect 59998 4060 60004 4072
rect 53800 4032 60004 4060
rect 53800 4020 53806 4032
rect 59998 4020 60004 4032
rect 60056 4020 60062 4072
rect 62022 4020 62028 4072
rect 62080 4060 62086 4072
rect 68646 4060 68652 4072
rect 62080 4032 68652 4060
rect 62080 4020 62086 4032
rect 68646 4020 68652 4032
rect 68704 4020 68710 4072
rect 69106 4020 69112 4072
rect 69164 4060 69170 4072
rect 76098 4060 76104 4072
rect 69164 4032 76104 4060
rect 69164 4020 69170 4032
rect 76098 4020 76104 4032
rect 76156 4020 76162 4072
rect 77386 4020 77392 4072
rect 77444 4060 77450 4072
rect 84378 4060 84384 4072
rect 77444 4032 84384 4060
rect 77444 4020 77450 4032
rect 84378 4020 84384 4032
rect 84436 4020 84442 4072
rect 125870 4020 125876 4072
rect 125928 4060 125934 4072
rect 133782 4060 133788 4072
rect 125928 4032 133788 4060
rect 125928 4020 125934 4032
rect 133782 4020 133788 4032
rect 133840 4020 133846 4072
rect 136450 4020 136456 4072
rect 136508 4060 136514 4072
rect 143442 4060 143448 4072
rect 136508 4032 143448 4060
rect 136508 4020 136514 4032
rect 143442 4020 143448 4032
rect 143500 4020 143506 4072
rect 155402 4020 155408 4072
rect 155460 4060 155466 4072
rect 161566 4060 161572 4072
rect 155460 4032 161572 4060
rect 155460 4020 155466 4032
rect 161566 4020 161572 4032
rect 161624 4020 161630 4072
rect 177850 4020 177856 4072
rect 177908 4060 177914 4072
rect 182174 4060 182180 4072
rect 177908 4032 182180 4060
rect 177908 4020 177914 4032
rect 182174 4020 182180 4032
rect 182232 4020 182238 4072
rect 187326 4020 187332 4072
rect 187384 4060 187390 4072
rect 190454 4060 190460 4072
rect 187384 4032 190460 4060
rect 187384 4020 187390 4032
rect 190454 4020 190460 4032
rect 190512 4020 190518 4072
rect 196802 4020 196808 4072
rect 196860 4060 196866 4072
rect 200206 4060 200212 4072
rect 196860 4032 200212 4060
rect 196860 4020 196866 4032
rect 200206 4020 200212 4032
rect 200264 4020 200270 4072
rect 340690 4020 340696 4072
rect 340748 4060 340754 4072
rect 345750 4060 345756 4072
rect 340748 4032 345756 4060
rect 340748 4020 340754 4032
rect 345750 4020 345756 4032
rect 345808 4020 345814 4072
rect 350442 4020 350448 4072
rect 350500 4060 350506 4072
rect 355226 4060 355232 4072
rect 350500 4032 355232 4060
rect 350500 4020 350506 4032
rect 355226 4020 355232 4032
rect 355284 4020 355290 4072
rect 361482 4020 361488 4072
rect 361540 4060 361546 4072
rect 367002 4060 367008 4072
rect 361540 4032 367008 4060
rect 361540 4020 361546 4032
rect 367002 4020 367008 4032
rect 367060 4020 367066 4072
rect 369762 4020 369768 4072
rect 369820 4060 369826 4072
rect 376478 4060 376484 4072
rect 369820 4032 376484 4060
rect 369820 4020 369826 4032
rect 376478 4020 376484 4032
rect 376536 4020 376542 4072
rect 406102 4020 406108 4072
rect 406160 4060 406166 4072
rect 415486 4060 415492 4072
rect 406160 4032 415492 4060
rect 406160 4020 406166 4032
rect 415486 4020 415492 4032
rect 415544 4020 415550 4072
rect 423030 4020 423036 4072
rect 423088 4060 423094 4072
rect 433242 4060 433248 4072
rect 423088 4032 433248 4060
rect 423088 4020 423094 4032
rect 433242 4020 433248 4032
rect 433300 4020 433306 4072
rect 524230 4020 524236 4072
rect 524288 4060 524294 4072
rect 529014 4060 529020 4072
rect 524288 4032 529020 4060
rect 524288 4020 524294 4032
rect 529014 4020 529020 4032
rect 529072 4020 529078 4072
rect 539410 4020 539416 4072
rect 539468 4060 539474 4072
rect 559742 4060 559748 4072
rect 539468 4032 559748 4060
rect 539468 4020 539474 4032
rect 559742 4020 559748 4032
rect 559800 4020 559806 4072
rect 9950 3952 9956 4004
rect 10008 3992 10014 4004
rect 22094 3992 22100 4004
rect 10008 3964 22100 3992
rect 10008 3952 10014 3964
rect 22094 3952 22100 3964
rect 22152 3952 22158 4004
rect 24210 3952 24216 4004
rect 24268 3992 24274 4004
rect 31662 3992 31668 4004
rect 24268 3964 31668 3992
rect 24268 3952 24274 3964
rect 31662 3952 31668 3964
rect 31720 3952 31726 4004
rect 54938 3952 54944 4004
rect 54996 3992 55002 4004
rect 60918 3992 60924 4004
rect 54996 3964 60924 3992
rect 54996 3952 55002 3964
rect 60918 3952 60924 3964
rect 60976 3952 60982 4004
rect 111610 3952 111616 4004
rect 111668 3992 111674 4004
rect 118050 3992 118056 4004
rect 111668 3964 118056 3992
rect 111668 3952 111674 3964
rect 118050 3952 118056 3964
rect 118108 3952 118114 4004
rect 118786 3952 118792 4004
rect 118844 3992 118850 4004
rect 126882 3992 126888 4004
rect 118844 3964 126888 3992
rect 118844 3952 118850 3964
rect 126882 3952 126888 3964
rect 126940 3952 126946 4004
rect 166074 3952 166080 4004
rect 166132 3992 166138 4004
rect 171134 3992 171140 4004
rect 166132 3964 171140 3992
rect 166132 3952 166138 3964
rect 171134 3952 171140 3964
rect 171192 3952 171198 4004
rect 313182 3952 313188 4004
rect 313240 3992 313246 4004
rect 316218 3992 316224 4004
rect 313240 3964 316224 3992
rect 313240 3952 313246 3964
rect 316218 3952 316224 3964
rect 316276 3952 316282 4004
rect 324130 3952 324136 4004
rect 324188 3992 324194 4004
rect 327994 3992 328000 4004
rect 324188 3964 328000 3992
rect 324188 3952 324194 3964
rect 327994 3952 328000 3964
rect 328052 3952 328058 4004
rect 360102 3952 360108 4004
rect 360160 3992 360166 4004
rect 365806 3992 365812 4004
rect 360160 3964 365812 3992
rect 360160 3952 360166 3964
rect 365806 3952 365812 3964
rect 365864 3952 365870 4004
rect 378042 3952 378048 4004
rect 378100 3992 378106 4004
rect 384758 3992 384764 4004
rect 378100 3964 384764 3992
rect 378100 3952 378106 3964
rect 384758 3952 384764 3964
rect 384816 3952 384822 4004
rect 389082 3952 389088 4004
rect 389140 3992 389146 4004
rect 396534 3992 396540 4004
rect 389140 3964 396540 3992
rect 389140 3952 389146 3964
rect 396534 3952 396540 3964
rect 396592 3952 396598 4004
rect 401502 3952 401508 4004
rect 401560 3992 401566 4004
rect 409598 3992 409604 4004
rect 401560 3964 409604 3992
rect 401560 3952 401566 3964
rect 409598 3952 409604 3964
rect 409656 3952 409662 4004
rect 412358 3952 412364 4004
rect 412416 3992 412422 4004
rect 421374 3992 421380 4004
rect 412416 3964 421380 3992
rect 412416 3952 412422 3964
rect 421374 3952 421380 3964
rect 421432 3952 421438 4004
rect 422294 3952 422300 4004
rect 422352 3992 422358 4004
rect 434438 3992 434444 4004
rect 422352 3964 434444 3992
rect 422352 3952 422358 3964
rect 434438 3952 434444 3964
rect 434496 3952 434502 4004
rect 488534 3952 488540 4004
rect 488592 3992 488598 4004
rect 491110 3992 491116 4004
rect 488592 3964 491116 3992
rect 488592 3952 488598 3964
rect 491110 3952 491116 3964
rect 491168 3952 491174 4004
rect 498194 3952 498200 4004
rect 498252 3992 498258 4004
rect 501782 3992 501788 4004
rect 498252 3964 501788 3992
rect 498252 3952 498258 3964
rect 501782 3952 501788 3964
rect 501840 3952 501846 4004
rect 533982 3952 533988 4004
rect 534040 3992 534046 4004
rect 538398 3992 538404 4004
rect 534040 3964 538404 3992
rect 534040 3952 534046 3964
rect 538398 3952 538404 3964
rect 538456 3952 538462 4004
rect 540514 3952 540520 4004
rect 540572 3992 540578 4004
rect 560846 3992 560852 4004
rect 540572 3964 560852 3992
rect 540572 3952 540578 3964
rect 560846 3952 560852 3964
rect 560904 3952 560910 4004
rect 4062 3884 4068 3936
rect 4120 3924 4126 3936
rect 16666 3924 16672 3936
rect 4120 3896 16672 3924
rect 4120 3884 4126 3896
rect 16666 3884 16672 3896
rect 16724 3884 16730 3936
rect 18046 3884 18052 3936
rect 18104 3924 18110 3936
rect 23658 3924 23664 3936
rect 18104 3896 23664 3924
rect 18104 3884 18110 3896
rect 23658 3884 23664 3896
rect 23716 3884 23722 3936
rect 44266 3884 44272 3936
rect 44324 3924 44330 3936
rect 52086 3924 52092 3936
rect 44324 3896 52092 3924
rect 44324 3884 44330 3896
rect 52086 3884 52092 3896
rect 52144 3884 52150 3936
rect 101030 3884 101036 3936
rect 101088 3924 101094 3936
rect 108206 3924 108212 3936
rect 101088 3896 108212 3924
rect 101088 3884 101094 3896
rect 108206 3884 108212 3896
rect 108264 3884 108270 3936
rect 332502 3884 332508 3936
rect 332560 3924 332566 3936
rect 336274 3924 336280 3936
rect 332560 3896 336280 3924
rect 332560 3884 332566 3896
rect 336274 3884 336280 3896
rect 336332 3884 336338 3936
rect 372614 3884 372620 3936
rect 372672 3924 372678 3936
rect 379974 3924 379980 3936
rect 372672 3896 379980 3924
rect 372672 3884 372678 3896
rect 379974 3884 379980 3896
rect 380032 3884 380038 3936
rect 392486 3884 392492 3936
rect 392544 3924 392550 3936
rect 401318 3924 401324 3936
rect 392544 3896 401324 3924
rect 392544 3884 392550 3896
rect 401318 3884 401324 3896
rect 401376 3884 401382 3936
rect 401410 3884 401416 3936
rect 401468 3924 401474 3936
rect 410794 3924 410800 3936
rect 401468 3896 410800 3924
rect 401468 3884 401474 3896
rect 410794 3884 410800 3896
rect 410852 3884 410858 3936
rect 411162 3884 411168 3936
rect 411220 3924 411226 3936
rect 420178 3924 420184 3936
rect 411220 3896 420184 3924
rect 411220 3884 411226 3896
rect 420178 3884 420184 3896
rect 420236 3884 420242 3936
rect 427722 3884 427728 3936
rect 427780 3924 427786 3936
rect 437934 3924 437940 3936
rect 427780 3896 437940 3924
rect 427780 3884 427786 3896
rect 437934 3884 437940 3896
rect 437992 3884 437998 3936
rect 534902 3884 534908 3936
rect 534960 3924 534966 3936
rect 539594 3924 539600 3936
rect 534960 3896 539600 3924
rect 534960 3884 534966 3896
rect 539594 3884 539600 3896
rect 539652 3884 539658 3936
rect 545022 3884 545028 3936
rect 545080 3924 545086 3936
rect 550266 3924 550272 3936
rect 545080 3896 550272 3924
rect 545080 3884 545086 3896
rect 550266 3884 550272 3896
rect 550324 3884 550330 3936
rect 552014 3884 552020 3936
rect 552072 3924 552078 3936
rect 553210 3924 553216 3936
rect 552072 3896 553216 3924
rect 552072 3884 552078 3896
rect 553210 3884 553216 3896
rect 553268 3884 553274 3936
rect 553394 3884 553400 3936
rect 553452 3924 553458 3936
rect 575106 3924 575112 3936
rect 553452 3896 575112 3924
rect 553452 3884 553458 3896
rect 575106 3884 575112 3896
rect 575164 3884 575170 3936
rect 2866 3816 2872 3868
rect 2924 3856 2930 3868
rect 17862 3856 17868 3868
rect 2924 3828 17868 3856
rect 2924 3816 2930 3828
rect 17862 3816 17868 3828
rect 17920 3816 17926 3868
rect 21818 3816 21824 3868
rect 21876 3856 21882 3868
rect 27614 3856 27620 3868
rect 21876 3828 27620 3856
rect 21876 3816 21882 3828
rect 27614 3816 27620 3828
rect 27672 3816 27678 3868
rect 31294 3816 31300 3868
rect 31352 3856 31358 3868
rect 37274 3856 37280 3868
rect 31352 3828 37280 3856
rect 31352 3816 31358 3828
rect 37274 3816 37280 3828
rect 37332 3816 37338 3868
rect 71498 3816 71504 3868
rect 71556 3856 71562 3868
rect 78582 3856 78588 3868
rect 71556 3828 78588 3856
rect 71556 3816 71562 3828
rect 78582 3816 78588 3828
rect 78640 3816 78646 3868
rect 80882 3816 80888 3868
rect 80940 3856 80946 3868
rect 87782 3856 87788 3868
rect 80940 3828 87788 3856
rect 80940 3816 80946 3828
rect 87782 3816 87788 3828
rect 87840 3816 87846 3868
rect 122282 3816 122288 3868
rect 122340 3856 122346 3868
rect 129642 3856 129648 3868
rect 122340 3828 129648 3856
rect 122340 3816 122346 3828
rect 129642 3816 129648 3828
rect 129700 3816 129706 3868
rect 141234 3816 141240 3868
rect 141292 3856 141298 3868
rect 147674 3856 147680 3868
rect 141292 3828 147680 3856
rect 141292 3816 141298 3828
rect 147674 3816 147680 3828
rect 147732 3816 147738 3868
rect 150618 3816 150624 3868
rect 150676 3856 150682 3868
rect 155954 3856 155960 3868
rect 150676 3828 155960 3856
rect 150676 3816 150682 3828
rect 155954 3816 155960 3828
rect 156012 3816 156018 3868
rect 167178 3816 167184 3868
rect 167236 3856 167242 3868
rect 172606 3856 172612 3868
rect 167236 3828 172612 3856
rect 167236 3816 167242 3828
rect 172606 3816 172612 3828
rect 172664 3816 172670 3868
rect 188522 3816 188528 3868
rect 188580 3856 188586 3868
rect 191926 3856 191932 3868
rect 188580 3828 191932 3856
rect 188580 3816 188586 3828
rect 191926 3816 191932 3828
rect 191984 3816 191990 3868
rect 286042 3816 286048 3868
rect 286100 3856 286106 3868
rect 287790 3856 287796 3868
rect 286100 3828 287796 3856
rect 286100 3816 286106 3828
rect 287790 3816 287796 3828
rect 287848 3816 287854 3868
rect 295518 3816 295524 3868
rect 295576 3856 295582 3868
rect 297266 3856 297272 3868
rect 295576 3828 297272 3856
rect 295576 3816 295582 3828
rect 297266 3816 297272 3828
rect 297324 3816 297330 3868
rect 305730 3816 305736 3868
rect 305788 3856 305794 3868
rect 307938 3856 307944 3868
rect 305788 3828 307944 3856
rect 305788 3816 305794 3828
rect 307938 3816 307944 3828
rect 307996 3816 308002 3868
rect 315850 3816 315856 3868
rect 315908 3856 315914 3868
rect 318518 3856 318524 3868
rect 315908 3828 318524 3856
rect 315908 3816 315914 3828
rect 318518 3816 318524 3828
rect 318576 3816 318582 3868
rect 362770 3816 362776 3868
rect 362828 3856 362834 3868
rect 368198 3856 368204 3868
rect 362828 3828 368204 3856
rect 362828 3816 362834 3828
rect 368198 3816 368204 3828
rect 368256 3816 368262 3868
rect 394786 3816 394792 3868
rect 394844 3856 394850 3868
rect 403618 3856 403624 3868
rect 394844 3828 403624 3856
rect 394844 3816 394850 3828
rect 403618 3816 403624 3828
rect 403676 3816 403682 3868
rect 407390 3816 407396 3868
rect 407448 3856 407454 3868
rect 417878 3856 417884 3868
rect 407448 3828 417884 3856
rect 407448 3816 407454 3828
rect 417878 3816 417884 3828
rect 417936 3816 417942 3868
rect 418062 3816 418068 3868
rect 418120 3856 418126 3868
rect 428458 3856 428464 3868
rect 418120 3828 428464 3856
rect 418120 3816 418126 3828
rect 428458 3816 428464 3828
rect 428516 3816 428522 3868
rect 429654 3816 429660 3868
rect 429712 3856 429718 3868
rect 441522 3856 441528 3868
rect 429712 3828 441528 3856
rect 429712 3816 429718 3828
rect 441522 3816 441528 3828
rect 441580 3816 441586 3868
rect 536006 3816 536012 3868
rect 536064 3856 536070 3868
rect 541986 3856 541992 3868
rect 536064 3828 541992 3856
rect 536064 3816 536070 3828
rect 541986 3816 541992 3828
rect 542044 3816 542050 3868
rect 542354 3816 542360 3868
rect 542412 3856 542418 3868
rect 549070 3856 549076 3868
rect 542412 3828 549076 3856
rect 542412 3816 542418 3828
rect 549070 3816 549076 3828
rect 549128 3816 549134 3868
rect 553486 3816 553492 3868
rect 553544 3856 553550 3868
rect 576302 3856 576308 3868
rect 553544 3828 576308 3856
rect 553544 3816 553550 3828
rect 576302 3816 576308 3828
rect 576360 3816 576366 3868
rect 566 3748 572 3800
rect 624 3788 630 3800
rect 13814 3788 13820 3800
rect 624 3760 13820 3788
rect 624 3748 630 3760
rect 13814 3748 13820 3760
rect 13872 3748 13878 3800
rect 15930 3748 15936 3800
rect 15988 3788 15994 3800
rect 23382 3788 23388 3800
rect 15988 3760 23388 3788
rect 15988 3748 15994 3760
rect 23382 3748 23388 3760
rect 23440 3748 23446 3800
rect 25314 3748 25320 3800
rect 25372 3788 25378 3800
rect 32766 3788 32772 3800
rect 25372 3760 32772 3788
rect 25372 3748 25378 3760
rect 32766 3748 32772 3760
rect 32824 3748 32830 3800
rect 34790 3748 34796 3800
rect 34848 3788 34854 3800
rect 41506 3788 41512 3800
rect 34848 3760 41512 3788
rect 34848 3748 34854 3760
rect 41506 3748 41512 3760
rect 41564 3748 41570 3800
rect 43070 3748 43076 3800
rect 43128 3788 43134 3800
rect 50982 3788 50988 3800
rect 43128 3760 50988 3788
rect 43128 3748 43134 3760
rect 50982 3748 50988 3760
rect 51040 3748 51046 3800
rect 51350 3748 51356 3800
rect 51408 3788 51414 3800
rect 59262 3788 59268 3800
rect 51408 3760 59268 3788
rect 51408 3748 51414 3760
rect 59262 3748 59268 3760
rect 59320 3748 59326 3800
rect 64322 3748 64328 3800
rect 64380 3788 64386 3800
rect 70946 3788 70952 3800
rect 64380 3760 70952 3788
rect 64380 3748 64386 3760
rect 70946 3748 70952 3760
rect 71004 3748 71010 3800
rect 99834 3748 99840 3800
rect 99892 3788 99898 3800
rect 106826 3788 106832 3800
rect 99892 3760 106832 3788
rect 99892 3748 99898 3760
rect 106826 3748 106832 3760
rect 106884 3748 106890 3800
rect 163682 3748 163688 3800
rect 163740 3788 163746 3800
rect 168374 3788 168380 3800
rect 163740 3760 168380 3788
rect 163740 3748 163746 3760
rect 168374 3748 168380 3760
rect 168432 3748 168438 3800
rect 335170 3748 335176 3800
rect 335228 3788 335234 3800
rect 338666 3788 338672 3800
rect 335228 3760 338672 3788
rect 335228 3748 335234 3760
rect 338666 3748 338672 3760
rect 338724 3748 338730 3800
rect 362862 3748 362868 3800
rect 362920 3788 362926 3800
rect 369394 3788 369400 3800
rect 362920 3760 369400 3788
rect 362920 3748 362926 3760
rect 369394 3748 369400 3760
rect 369452 3748 369458 3800
rect 372154 3748 372160 3800
rect 372212 3788 372218 3800
rect 378870 3788 378876 3800
rect 372212 3760 378876 3788
rect 372212 3748 372218 3760
rect 378870 3748 378876 3760
rect 378928 3748 378934 3800
rect 379422 3748 379428 3800
rect 379480 3788 379486 3800
rect 387150 3788 387156 3800
rect 379480 3760 387156 3788
rect 379480 3748 379486 3760
rect 387150 3748 387156 3760
rect 387208 3748 387214 3800
rect 391842 3748 391848 3800
rect 391900 3788 391906 3800
rect 400030 3788 400036 3800
rect 391900 3760 400036 3788
rect 391900 3748 391906 3760
rect 400030 3748 400036 3760
rect 400088 3748 400094 3800
rect 400122 3748 400128 3800
rect 400180 3788 400186 3800
rect 408402 3788 408408 3800
rect 400180 3760 408408 3788
rect 400180 3748 400186 3760
rect 408402 3748 408408 3760
rect 408460 3748 408466 3800
rect 420822 3748 420828 3800
rect 420880 3788 420886 3800
rect 430850 3788 430856 3800
rect 420880 3760 430856 3788
rect 420880 3748 420886 3760
rect 430850 3748 430856 3760
rect 430908 3748 430914 3800
rect 430942 3748 430948 3800
rect 431000 3788 431006 3800
rect 442626 3788 442632 3800
rect 431000 3760 442632 3788
rect 431000 3748 431006 3760
rect 442626 3748 442632 3760
rect 442684 3748 442690 3800
rect 478874 3748 478880 3800
rect 478932 3788 478938 3800
rect 481726 3788 481732 3800
rect 478932 3760 481732 3788
rect 478932 3748 478938 3760
rect 481726 3748 481732 3760
rect 481784 3748 481790 3800
rect 538030 3748 538036 3800
rect 538088 3788 538094 3800
rect 543182 3788 543188 3800
rect 538088 3760 543188 3788
rect 538088 3748 538094 3760
rect 543182 3748 543188 3760
rect 543240 3748 543246 3800
rect 550634 3748 550640 3800
rect 550692 3788 550698 3800
rect 552750 3788 552756 3800
rect 550692 3760 552756 3788
rect 550692 3748 550698 3760
rect 552750 3748 552756 3760
rect 552808 3748 552814 3800
rect 554774 3748 554780 3800
rect 554832 3788 554838 3800
rect 577406 3788 577412 3800
rect 554832 3760 577412 3788
rect 554832 3748 554838 3760
rect 577406 3748 577412 3760
rect 577464 3748 577470 3800
rect 11146 3680 11152 3732
rect 11204 3720 11210 3732
rect 26234 3720 26240 3732
rect 11204 3692 26240 3720
rect 11204 3680 11210 3692
rect 26234 3680 26240 3692
rect 26292 3680 26298 3732
rect 32398 3680 32404 3732
rect 32456 3720 32462 3732
rect 39298 3720 39304 3732
rect 32456 3692 39304 3720
rect 32456 3680 32462 3692
rect 39298 3680 39304 3692
rect 39356 3680 39362 3732
rect 41874 3680 41880 3732
rect 41932 3720 41938 3732
rect 49602 3720 49608 3732
rect 41932 3692 49608 3720
rect 41932 3680 41938 3692
rect 49602 3680 49608 3692
rect 49660 3680 49666 3732
rect 73798 3680 73804 3732
rect 73856 3720 73862 3732
rect 80514 3720 80520 3732
rect 73856 3692 80520 3720
rect 73856 3680 73862 3692
rect 80514 3680 80520 3692
rect 80572 3680 80578 3732
rect 92750 3680 92756 3732
rect 92808 3720 92814 3732
rect 99466 3720 99472 3732
rect 92808 3692 99472 3720
rect 92808 3680 92814 3692
rect 99466 3680 99472 3692
rect 99524 3680 99530 3732
rect 106918 3680 106924 3732
rect 106976 3720 106982 3732
rect 113266 3720 113272 3732
rect 106976 3692 113272 3720
rect 106976 3680 106982 3692
rect 113266 3680 113272 3692
rect 113324 3680 113330 3732
rect 121086 3680 121092 3732
rect 121144 3720 121150 3732
rect 128262 3720 128268 3732
rect 121144 3692 128268 3720
rect 121144 3680 121150 3692
rect 128262 3680 128268 3692
rect 128320 3680 128326 3732
rect 140038 3680 140044 3732
rect 140096 3720 140102 3732
rect 146294 3720 146300 3732
rect 140096 3692 146300 3720
rect 140096 3680 140102 3692
rect 146294 3680 146300 3692
rect 146352 3680 146358 3732
rect 148318 3680 148324 3732
rect 148376 3720 148382 3732
rect 154574 3720 154580 3732
rect 148376 3692 154580 3720
rect 148376 3680 148382 3692
rect 154574 3680 154580 3692
rect 154632 3680 154638 3732
rect 160094 3680 160100 3732
rect 160152 3720 160158 3732
rect 165614 3720 165620 3732
rect 160152 3692 165620 3720
rect 160152 3680 160158 3692
rect 165614 3680 165620 3692
rect 165672 3680 165678 3732
rect 171962 3680 171968 3732
rect 172020 3720 172026 3732
rect 176654 3720 176660 3732
rect 172020 3692 176660 3720
rect 172020 3680 172026 3692
rect 176654 3680 176660 3692
rect 176712 3680 176718 3732
rect 304442 3680 304448 3732
rect 304500 3720 304506 3732
rect 306742 3720 306748 3732
rect 304500 3692 306748 3720
rect 304500 3680 304506 3692
rect 306742 3680 306748 3692
rect 306800 3680 306806 3732
rect 354490 3680 354496 3732
rect 354548 3720 354554 3732
rect 359918 3720 359924 3732
rect 354548 3692 359924 3720
rect 354548 3680 354554 3692
rect 359918 3680 359924 3692
rect 359976 3680 359982 3732
rect 382918 3680 382924 3732
rect 382976 3720 382982 3732
rect 390646 3720 390652 3732
rect 382976 3692 390652 3720
rect 382976 3680 382982 3692
rect 390646 3680 390652 3692
rect 390704 3680 390710 3732
rect 394878 3680 394884 3732
rect 394936 3720 394942 3732
rect 404814 3720 404820 3732
rect 394936 3692 404820 3720
rect 394936 3680 394942 3692
rect 404814 3680 404820 3692
rect 404872 3680 404878 3732
rect 407022 3680 407028 3732
rect 407080 3720 407086 3732
rect 416682 3720 416688 3732
rect 407080 3692 416688 3720
rect 407080 3680 407086 3692
rect 416682 3680 416688 3692
rect 416740 3680 416746 3732
rect 423766 3680 423772 3732
rect 423824 3720 423830 3732
rect 435542 3720 435548 3732
rect 423824 3692 435548 3720
rect 423824 3680 423830 3692
rect 435542 3680 435548 3692
rect 435600 3680 435606 3732
rect 438670 3680 438676 3732
rect 438728 3720 438734 3732
rect 449802 3720 449808 3732
rect 438728 3692 449808 3720
rect 438728 3680 438734 3692
rect 449802 3680 449808 3692
rect 449860 3680 449866 3732
rect 527910 3680 527916 3732
rect 527968 3720 527974 3732
rect 532510 3720 532516 3732
rect 527968 3692 532516 3720
rect 527968 3680 527974 3692
rect 532510 3680 532516 3692
rect 532568 3680 532574 3732
rect 545758 3680 545764 3732
rect 545816 3720 545822 3732
rect 551462 3720 551468 3732
rect 545816 3692 551468 3720
rect 545816 3680 545822 3692
rect 551462 3680 551468 3692
rect 551520 3680 551526 3732
rect 556154 3680 556160 3732
rect 556212 3720 556218 3732
rect 578602 3720 578608 3732
rect 556212 3692 578608 3720
rect 556212 3680 556218 3692
rect 578602 3680 578608 3692
rect 578660 3680 578666 3732
rect 6454 3612 6460 3664
rect 6512 3652 6518 3664
rect 22186 3652 22192 3664
rect 6512 3624 22192 3652
rect 6512 3612 6518 3624
rect 22186 3612 22192 3624
rect 22244 3612 22250 3664
rect 23014 3612 23020 3664
rect 23072 3652 23078 3664
rect 29914 3652 29920 3664
rect 23072 3624 29920 3652
rect 23072 3612 23078 3624
rect 29914 3612 29920 3624
rect 29972 3612 29978 3664
rect 63218 3612 63224 3664
rect 63276 3652 63282 3664
rect 69934 3652 69940 3664
rect 63276 3624 69940 3652
rect 63276 3612 63282 3624
rect 69934 3612 69940 3624
rect 69992 3612 69998 3664
rect 72602 3612 72608 3664
rect 72660 3652 72666 3664
rect 79962 3652 79968 3664
rect 72660 3624 79968 3652
rect 72660 3612 72666 3624
rect 79962 3612 79968 3624
rect 80020 3612 80026 3664
rect 104526 3612 104532 3664
rect 104584 3652 104590 3664
rect 110506 3652 110512 3664
rect 104584 3624 110512 3652
rect 104584 3612 104590 3624
rect 110506 3612 110512 3624
rect 110564 3612 110570 3664
rect 130562 3612 130568 3664
rect 130620 3652 130626 3664
rect 137922 3652 137928 3664
rect 130620 3624 137928 3652
rect 130620 3612 130626 3624
rect 137922 3612 137928 3624
rect 137980 3612 137986 3664
rect 138842 3612 138848 3664
rect 138900 3652 138906 3664
rect 145098 3652 145104 3664
rect 138900 3624 145104 3652
rect 138900 3612 138906 3624
rect 145098 3612 145104 3624
rect 145156 3612 145162 3664
rect 158898 3612 158904 3664
rect 158956 3652 158962 3664
rect 164234 3652 164240 3664
rect 158956 3624 164240 3652
rect 158956 3612 158962 3624
rect 164234 3612 164240 3624
rect 164292 3612 164298 3664
rect 169570 3612 169576 3664
rect 169628 3652 169634 3664
rect 173894 3652 173900 3664
rect 169628 3624 173900 3652
rect 169628 3612 169634 3624
rect 173894 3612 173900 3624
rect 173952 3612 173958 3664
rect 353202 3612 353208 3664
rect 353260 3652 353266 3664
rect 358722 3652 358728 3664
rect 353260 3624 358728 3652
rect 353260 3612 353266 3624
rect 358722 3612 358728 3624
rect 358780 3612 358786 3664
rect 363322 3612 363328 3664
rect 363380 3652 363386 3664
rect 370590 3652 370596 3664
rect 363380 3624 370596 3652
rect 363380 3612 363386 3624
rect 370590 3612 370596 3624
rect 370648 3612 370654 3664
rect 371142 3612 371148 3664
rect 371200 3652 371206 3664
rect 377674 3652 377680 3664
rect 371200 3624 377680 3652
rect 371200 3612 371206 3624
rect 377674 3612 377680 3624
rect 377732 3612 377738 3664
rect 385034 3612 385040 3664
rect 385092 3652 385098 3664
rect 385092 3624 388484 3652
rect 385092 3612 385098 3624
rect 12342 3544 12348 3596
rect 12400 3584 12406 3596
rect 27798 3584 27804 3596
rect 12400 3556 27804 3584
rect 12400 3544 12406 3556
rect 27798 3544 27804 3556
rect 27856 3544 27862 3596
rect 33594 3544 33600 3596
rect 33652 3584 33658 3596
rect 41322 3584 41328 3596
rect 33652 3556 41328 3584
rect 33652 3544 33658 3556
rect 41322 3544 41328 3556
rect 41380 3544 41386 3596
rect 59630 3544 59636 3596
rect 59688 3584 59694 3596
rect 66346 3584 66352 3596
rect 59688 3556 66352 3584
rect 59688 3544 59694 3556
rect 66346 3544 66352 3556
rect 66404 3544 66410 3596
rect 82078 3544 82084 3596
rect 82136 3584 82142 3596
rect 89622 3584 89628 3596
rect 82136 3556 89628 3584
rect 82136 3544 82142 3556
rect 89622 3544 89628 3556
rect 89680 3544 89686 3596
rect 90358 3544 90364 3596
rect 90416 3584 90422 3596
rect 97166 3584 97172 3596
rect 90416 3556 97172 3584
rect 90416 3544 90422 3556
rect 97166 3544 97172 3556
rect 97224 3544 97230 3596
rect 109310 3544 109316 3596
rect 109368 3584 109374 3596
rect 117222 3584 117228 3596
rect 109368 3556 117228 3584
rect 109368 3544 109374 3556
rect 117222 3544 117228 3556
rect 117280 3544 117286 3596
rect 131758 3544 131764 3596
rect 131816 3584 131822 3596
rect 139302 3584 139308 3596
rect 131816 3556 139308 3584
rect 131816 3544 131822 3556
rect 139302 3544 139308 3556
rect 139360 3544 139366 3596
rect 170766 3544 170772 3596
rect 170824 3584 170830 3596
rect 175274 3584 175280 3596
rect 170824 3556 175280 3584
rect 170824 3544 170830 3556
rect 175274 3544 175280 3556
rect 175332 3544 175338 3596
rect 180242 3544 180248 3596
rect 180300 3584 180306 3596
rect 183646 3584 183652 3596
rect 180300 3556 183652 3584
rect 180300 3544 180306 3556
rect 183646 3544 183652 3556
rect 183704 3544 183710 3596
rect 259454 3544 259460 3596
rect 259512 3584 259518 3596
rect 260650 3584 260656 3596
rect 259512 3556 260656 3584
rect 259512 3544 259518 3556
rect 260650 3544 260656 3556
rect 260708 3544 260714 3596
rect 303154 3544 303160 3596
rect 303212 3584 303218 3596
rect 305546 3584 305552 3596
rect 303212 3556 305552 3584
rect 303212 3544 303218 3556
rect 305546 3544 305552 3556
rect 305604 3544 305610 3596
rect 346394 3544 346400 3596
rect 346452 3584 346458 3596
rect 352834 3584 352840 3596
rect 346452 3556 352840 3584
rect 346452 3544 346458 3556
rect 352834 3544 352840 3556
rect 352892 3544 352898 3596
rect 368382 3544 368388 3596
rect 368440 3584 368446 3596
rect 374086 3584 374092 3596
rect 368440 3556 374092 3584
rect 368440 3544 368446 3556
rect 374086 3544 374092 3556
rect 374144 3544 374150 3596
rect 380802 3544 380808 3596
rect 380860 3584 380866 3596
rect 388254 3584 388260 3596
rect 380860 3556 388260 3584
rect 380860 3544 380866 3556
rect 388254 3544 388260 3556
rect 388312 3544 388318 3596
rect 388456 3584 388484 3624
rect 402882 3612 402888 3664
rect 402940 3652 402946 3664
rect 411898 3652 411904 3664
rect 402940 3624 411904 3652
rect 402940 3612 402946 3624
rect 411898 3612 411904 3624
rect 411956 3612 411962 3664
rect 412542 3612 412548 3664
rect 412600 3652 412606 3664
rect 422570 3652 422576 3664
rect 412600 3624 422576 3652
rect 412600 3612 412606 3624
rect 422570 3612 422576 3624
rect 422628 3612 422634 3664
rect 427814 3612 427820 3664
rect 427872 3652 427878 3664
rect 439130 3652 439136 3664
rect 427872 3624 439136 3652
rect 427872 3612 427878 3624
rect 439130 3612 439136 3624
rect 439188 3612 439194 3664
rect 551830 3612 551836 3664
rect 551888 3652 551894 3664
rect 558546 3652 558552 3664
rect 551888 3624 558552 3652
rect 551888 3612 551894 3624
rect 558546 3612 558552 3624
rect 558604 3612 558610 3664
rect 560294 3612 560300 3664
rect 560352 3652 560358 3664
rect 583386 3652 583392 3664
rect 560352 3624 583392 3652
rect 560352 3612 560358 3624
rect 583386 3612 583392 3624
rect 583444 3612 583450 3664
rect 394234 3584 394240 3596
rect 388456 3556 394240 3584
rect 394234 3544 394240 3556
rect 394292 3544 394298 3596
rect 396258 3544 396264 3596
rect 396316 3584 396322 3596
rect 396316 3556 402974 3584
rect 396316 3544 396322 3556
rect 7650 3476 7656 3528
rect 7708 3516 7714 3528
rect 18046 3516 18052 3528
rect 7708 3488 18052 3516
rect 7708 3476 7714 3488
rect 18046 3476 18052 3488
rect 18104 3476 18110 3528
rect 18230 3476 18236 3528
rect 18288 3516 18294 3528
rect 25038 3516 25044 3528
rect 18288 3488 25044 3516
rect 18288 3476 18294 3488
rect 25038 3476 25044 3488
rect 25096 3476 25102 3528
rect 26510 3476 26516 3528
rect 26568 3516 26574 3528
rect 33778 3516 33784 3528
rect 26568 3488 33784 3516
rect 26568 3476 26574 3488
rect 33778 3476 33784 3488
rect 33836 3476 33842 3528
rect 37182 3476 37188 3528
rect 37240 3516 37246 3528
rect 43438 3516 43444 3528
rect 37240 3488 43444 3516
rect 37240 3476 37246 3488
rect 43438 3476 43444 3488
rect 43496 3476 43502 3528
rect 47854 3476 47860 3528
rect 47912 3516 47918 3528
rect 53926 3516 53932 3528
rect 47912 3488 53932 3516
rect 47912 3476 47918 3488
rect 53926 3476 53932 3488
rect 53984 3476 53990 3528
rect 57238 3476 57244 3528
rect 57296 3516 57302 3528
rect 63494 3516 63500 3528
rect 57296 3488 63500 3516
rect 57296 3476 57302 3488
rect 63494 3476 63500 3488
rect 63552 3476 63558 3528
rect 74994 3476 75000 3528
rect 75052 3516 75058 3528
rect 81526 3516 81532 3528
rect 75052 3488 81532 3516
rect 75052 3476 75058 3488
rect 81526 3476 81532 3488
rect 81584 3476 81590 3528
rect 83274 3476 83280 3528
rect 83332 3516 83338 3528
rect 90174 3516 90180 3528
rect 83332 3488 90180 3516
rect 83332 3476 83338 3488
rect 90174 3476 90180 3488
rect 90232 3476 90238 3528
rect 91554 3476 91560 3528
rect 91612 3516 91618 3528
rect 98454 3516 98460 3528
rect 91612 3488 98460 3516
rect 91612 3476 91618 3488
rect 98454 3476 98460 3488
rect 98512 3476 98518 3528
rect 103330 3476 103336 3528
rect 103388 3516 103394 3528
rect 109126 3516 109132 3528
rect 103388 3488 109132 3516
rect 103388 3476 103394 3488
rect 109126 3476 109132 3488
rect 109184 3476 109190 3528
rect 112806 3476 112812 3528
rect 112864 3516 112870 3528
rect 118694 3516 118700 3528
rect 112864 3488 118700 3516
rect 112864 3476 112870 3488
rect 118694 3476 118700 3488
rect 118752 3476 118758 3528
rect 151814 3476 151820 3528
rect 151872 3516 151878 3528
rect 157334 3516 157340 3528
rect 151872 3488 157340 3516
rect 151872 3476 151878 3488
rect 157334 3476 157340 3488
rect 157392 3476 157398 3528
rect 168374 3476 168380 3528
rect 168432 3516 168438 3528
rect 172514 3516 172520 3528
rect 168432 3488 172520 3516
rect 168432 3476 168438 3488
rect 172514 3476 172520 3488
rect 172572 3476 172578 3528
rect 174262 3476 174268 3528
rect 174320 3516 174326 3528
rect 178126 3516 178132 3528
rect 174320 3488 178132 3516
rect 174320 3476 174326 3488
rect 178126 3476 178132 3488
rect 178184 3476 178190 3528
rect 179046 3476 179052 3528
rect 179104 3516 179110 3528
rect 183554 3516 183560 3528
rect 179104 3488 183560 3516
rect 179104 3476 179110 3488
rect 183554 3476 183560 3488
rect 183612 3476 183618 3528
rect 183738 3476 183744 3528
rect 183796 3516 183802 3528
rect 187694 3516 187700 3528
rect 183796 3488 187700 3516
rect 183796 3476 183802 3488
rect 187694 3476 187700 3488
rect 187752 3476 187758 3528
rect 189718 3476 189724 3528
rect 189776 3516 189782 3528
rect 193306 3516 193312 3528
rect 189776 3488 193312 3516
rect 189776 3476 189782 3488
rect 193306 3476 193312 3488
rect 193364 3476 193370 3528
rect 291010 3476 291016 3528
rect 291068 3516 291074 3528
rect 292574 3516 292580 3528
rect 291068 3488 292580 3516
rect 291068 3476 291074 3488
rect 292574 3476 292580 3488
rect 292632 3476 292638 3528
rect 292942 3476 292948 3528
rect 293000 3516 293006 3528
rect 294874 3516 294880 3528
rect 293000 3488 294880 3516
rect 293000 3476 293006 3488
rect 294874 3476 294880 3488
rect 294932 3476 294938 3528
rect 300670 3476 300676 3528
rect 300728 3516 300734 3528
rect 301958 3516 301964 3528
rect 300728 3488 301964 3516
rect 300728 3476 300734 3488
rect 301958 3476 301964 3488
rect 302016 3476 302022 3528
rect 306926 3476 306932 3528
rect 306984 3516 306990 3528
rect 309042 3516 309048 3528
rect 306984 3488 309048 3516
rect 306984 3476 306990 3488
rect 309042 3476 309048 3488
rect 309100 3476 309106 3528
rect 310422 3476 310428 3528
rect 310480 3516 310486 3528
rect 312630 3516 312636 3528
rect 310480 3488 312636 3516
rect 310480 3476 310486 3488
rect 312630 3476 312636 3488
rect 312688 3476 312694 3528
rect 316034 3476 316040 3528
rect 316092 3516 316098 3528
rect 319714 3516 319720 3528
rect 316092 3488 319720 3516
rect 316092 3476 316098 3488
rect 319714 3476 319720 3488
rect 319772 3476 319778 3528
rect 322842 3476 322848 3528
rect 322900 3516 322906 3528
rect 325602 3516 325608 3528
rect 322900 3488 325608 3516
rect 322900 3476 322906 3488
rect 325602 3476 325608 3488
rect 325660 3476 325666 3528
rect 329742 3476 329748 3528
rect 329800 3516 329806 3528
rect 332686 3516 332692 3528
rect 329800 3488 332692 3516
rect 329800 3476 329806 3488
rect 332686 3476 332692 3488
rect 332744 3476 332750 3528
rect 334250 3476 334256 3528
rect 334308 3516 334314 3528
rect 339862 3516 339868 3528
rect 334308 3488 339868 3516
rect 334308 3476 334314 3488
rect 339862 3476 339868 3488
rect 339920 3476 339926 3528
rect 343542 3476 343548 3528
rect 343600 3516 343606 3528
rect 348050 3516 348056 3528
rect 343600 3488 348056 3516
rect 343600 3476 343606 3488
rect 348050 3476 348056 3488
rect 348108 3476 348114 3528
rect 355042 3476 355048 3528
rect 355100 3516 355106 3528
rect 361114 3516 361120 3528
rect 355100 3488 361120 3516
rect 355100 3476 355106 3488
rect 361114 3476 361120 3488
rect 361172 3476 361178 3528
rect 390462 3476 390468 3528
rect 390520 3516 390526 3528
rect 398926 3516 398932 3528
rect 390520 3488 398932 3516
rect 390520 3476 390526 3488
rect 398926 3476 398932 3488
rect 398984 3476 398990 3528
rect 402946 3516 402974 3556
rect 403434 3544 403440 3596
rect 403492 3584 403498 3596
rect 413094 3584 413100 3596
rect 403492 3556 413100 3584
rect 403492 3544 403498 3556
rect 413094 3544 413100 3556
rect 413152 3544 413158 3596
rect 420914 3544 420920 3596
rect 420972 3584 420978 3596
rect 432046 3584 432052 3596
rect 420972 3556 432052 3584
rect 420972 3544 420978 3556
rect 432046 3544 432052 3556
rect 432104 3544 432110 3596
rect 432230 3544 432236 3596
rect 432288 3584 432294 3596
rect 443822 3584 443828 3596
rect 432288 3556 443828 3584
rect 432288 3544 432294 3556
rect 443822 3544 443828 3556
rect 443880 3544 443886 3596
rect 471974 3544 471980 3596
rect 472032 3584 472038 3596
rect 473446 3584 473452 3596
rect 472032 3556 473452 3584
rect 472032 3544 472038 3556
rect 473446 3544 473452 3556
rect 473504 3544 473510 3596
rect 491386 3544 491392 3596
rect 491444 3584 491450 3596
rect 494698 3584 494704 3596
rect 491444 3556 494704 3584
rect 491444 3544 491450 3556
rect 494698 3544 494704 3556
rect 494756 3544 494762 3596
rect 507854 3544 507860 3596
rect 507912 3584 507918 3596
rect 512454 3584 512460 3596
rect 507912 3556 512460 3584
rect 507912 3544 507918 3556
rect 512454 3544 512460 3556
rect 512512 3544 512518 3596
rect 516042 3544 516048 3596
rect 516100 3584 516106 3596
rect 519538 3584 519544 3596
rect 516100 3556 519544 3584
rect 516100 3544 516106 3556
rect 519538 3544 519544 3556
rect 519596 3544 519602 3596
rect 526438 3544 526444 3596
rect 526496 3584 526502 3596
rect 531314 3584 531320 3596
rect 526496 3556 531320 3584
rect 526496 3544 526502 3556
rect 531314 3544 531320 3556
rect 531372 3544 531378 3596
rect 531406 3544 531412 3596
rect 531464 3584 531470 3596
rect 531464 3556 534074 3584
rect 531464 3544 531470 3556
rect 406010 3516 406016 3528
rect 402946 3488 406016 3516
rect 406010 3476 406016 3488
rect 406068 3476 406074 3528
rect 412634 3476 412640 3528
rect 412692 3516 412698 3528
rect 423766 3516 423772 3528
rect 412692 3488 423772 3516
rect 412692 3476 412698 3488
rect 423766 3476 423772 3488
rect 423824 3476 423830 3528
rect 426066 3476 426072 3528
rect 426124 3516 426130 3528
rect 436738 3516 436744 3528
rect 426124 3488 436744 3516
rect 426124 3476 426130 3488
rect 436738 3476 436744 3488
rect 436796 3476 436802 3528
rect 438854 3476 438860 3528
rect 438912 3516 438918 3528
rect 450906 3516 450912 3528
rect 438912 3488 450912 3516
rect 438912 3476 438918 3488
rect 450906 3476 450912 3488
rect 450964 3476 450970 3528
rect 462314 3476 462320 3528
rect 462372 3516 462378 3528
rect 463970 3516 463976 3528
rect 462372 3488 463976 3516
rect 462372 3476 462378 3488
rect 463970 3476 463976 3488
rect 464028 3476 464034 3528
rect 467834 3476 467840 3528
rect 467892 3516 467898 3528
rect 469858 3516 469864 3528
rect 467892 3488 469864 3516
rect 467892 3476 467898 3488
rect 469858 3476 469864 3488
rect 469916 3476 469922 3528
rect 474642 3476 474648 3528
rect 474700 3516 474706 3528
rect 475746 3516 475752 3528
rect 474700 3488 475752 3516
rect 474700 3476 474706 3488
rect 475746 3476 475752 3488
rect 475804 3476 475810 3528
rect 476298 3476 476304 3528
rect 476356 3516 476362 3528
rect 478138 3516 478144 3528
rect 476356 3488 478144 3516
rect 476356 3476 476362 3488
rect 478138 3476 478144 3488
rect 478196 3476 478202 3528
rect 480622 3476 480628 3528
rect 480680 3516 480686 3528
rect 482830 3516 482836 3528
rect 480680 3488 482836 3516
rect 480680 3476 480686 3488
rect 482830 3476 482836 3488
rect 482888 3476 482894 3528
rect 484302 3476 484308 3528
rect 484360 3516 484366 3528
rect 485222 3516 485228 3528
rect 484360 3488 485228 3516
rect 484360 3476 484366 3488
rect 485222 3476 485228 3488
rect 485280 3476 485286 3528
rect 490098 3476 490104 3528
rect 490156 3516 490162 3528
rect 492306 3516 492312 3528
rect 490156 3488 492312 3516
rect 490156 3476 490162 3488
rect 492306 3476 492312 3488
rect 492364 3476 492370 3528
rect 496446 3476 496452 3528
rect 496504 3516 496510 3528
rect 499390 3516 499396 3528
rect 496504 3488 499396 3516
rect 496504 3476 496510 3488
rect 499390 3476 499396 3488
rect 499448 3476 499454 3528
rect 499666 3476 499672 3528
rect 499724 3516 499730 3528
rect 502978 3516 502984 3528
rect 499724 3488 502984 3516
rect 499724 3476 499730 3488
rect 502978 3476 502984 3488
rect 503036 3476 503042 3528
rect 505554 3476 505560 3528
rect 505612 3516 505618 3528
rect 508866 3516 508872 3528
rect 505612 3488 508872 3516
rect 505612 3476 505618 3488
rect 508866 3476 508872 3488
rect 508924 3476 508930 3528
rect 513282 3476 513288 3528
rect 513340 3516 513346 3528
rect 515950 3516 515956 3528
rect 513340 3488 515956 3516
rect 513340 3476 513346 3488
rect 515950 3476 515956 3488
rect 516008 3476 516014 3528
rect 517514 3476 517520 3528
rect 517572 3516 517578 3528
rect 521838 3516 521844 3528
rect 517572 3488 521844 3516
rect 517572 3476 517578 3488
rect 521838 3476 521844 3488
rect 521896 3476 521902 3528
rect 524322 3476 524328 3528
rect 524380 3516 524386 3528
rect 527818 3516 527824 3528
rect 524380 3488 527824 3516
rect 524380 3476 524386 3488
rect 527818 3476 527824 3488
rect 527876 3476 527882 3528
rect 528554 3476 528560 3528
rect 528612 3516 528618 3528
rect 533706 3516 533712 3528
rect 528612 3488 533712 3516
rect 528612 3476 528618 3488
rect 533706 3476 533712 3488
rect 533764 3476 533770 3528
rect 534046 3516 534074 3556
rect 538858 3544 538864 3596
rect 538916 3584 538922 3596
rect 544378 3584 544384 3596
rect 538916 3556 544384 3584
rect 538916 3544 538922 3556
rect 544378 3544 544384 3556
rect 544436 3544 544442 3596
rect 547874 3544 547880 3596
rect 547932 3584 547938 3596
rect 554958 3584 554964 3596
rect 547932 3556 554964 3584
rect 547932 3544 547938 3556
rect 554958 3544 554964 3556
rect 555016 3544 555022 3596
rect 558914 3544 558920 3596
rect 558972 3584 558978 3596
rect 580994 3584 581000 3596
rect 558972 3556 581000 3584
rect 558972 3544 558978 3556
rect 580994 3544 581000 3556
rect 581052 3544 581058 3596
rect 534046 3488 543734 3516
rect 1670 3408 1676 3460
rect 1728 3448 1734 3460
rect 18138 3448 18144 3460
rect 1728 3420 18144 3448
rect 1728 3408 1734 3420
rect 18138 3408 18144 3420
rect 18196 3408 18202 3460
rect 19426 3408 19432 3460
rect 19484 3448 19490 3460
rect 26418 3448 26424 3460
rect 19484 3420 26424 3448
rect 19484 3408 19490 3420
rect 26418 3408 26424 3420
rect 26476 3408 26482 3460
rect 45462 3408 45468 3460
rect 45520 3448 45526 3460
rect 52270 3448 52276 3460
rect 45520 3420 52276 3448
rect 45520 3408 45526 3420
rect 52270 3408 52276 3420
rect 52328 3408 52334 3460
rect 52546 3408 52552 3460
rect 52604 3448 52610 3460
rect 60550 3448 60556 3460
rect 52604 3420 60556 3448
rect 52604 3408 52610 3420
rect 60550 3408 60556 3420
rect 60608 3408 60614 3460
rect 60826 3408 60832 3460
rect 60884 3448 60890 3460
rect 68922 3448 68928 3460
rect 60884 3420 68928 3448
rect 60884 3408 60890 3420
rect 68922 3408 68928 3420
rect 68980 3408 68986 3460
rect 70302 3408 70308 3460
rect 70360 3448 70366 3460
rect 75914 3448 75920 3460
rect 70360 3420 75920 3448
rect 70360 3408 70366 3420
rect 75914 3408 75920 3420
rect 75972 3408 75978 3460
rect 85666 3408 85672 3460
rect 85724 3448 85730 3460
rect 92566 3448 92572 3460
rect 85724 3420 92572 3448
rect 85724 3408 85730 3420
rect 92566 3408 92572 3420
rect 92624 3408 92630 3460
rect 95142 3408 95148 3460
rect 95200 3448 95206 3460
rect 100846 3448 100852 3460
rect 95200 3420 100852 3448
rect 95200 3408 95206 3420
rect 100846 3408 100852 3420
rect 100904 3408 100910 3460
rect 102226 3408 102232 3460
rect 102284 3448 102290 3460
rect 109218 3448 109224 3460
rect 102284 3420 109224 3448
rect 102284 3408 102290 3420
rect 109218 3408 109224 3420
rect 109276 3408 109282 3460
rect 110506 3408 110512 3460
rect 110564 3448 110570 3460
rect 118602 3448 118608 3460
rect 110564 3420 118608 3448
rect 110564 3408 110570 3420
rect 118602 3408 118608 3420
rect 118660 3408 118666 3460
rect 119890 3408 119896 3460
rect 119948 3448 119954 3460
rect 126514 3448 126520 3460
rect 119948 3420 126520 3448
rect 119948 3408 119954 3420
rect 126514 3408 126520 3420
rect 126572 3408 126578 3460
rect 129366 3408 129372 3460
rect 129424 3448 129430 3460
rect 136542 3448 136548 3460
rect 129424 3420 136548 3448
rect 129424 3408 129430 3420
rect 136542 3408 136548 3420
rect 136600 3408 136606 3460
rect 142430 3408 142436 3460
rect 142488 3448 142494 3460
rect 149054 3448 149060 3460
rect 142488 3420 149060 3448
rect 142488 3408 142494 3420
rect 149054 3408 149060 3420
rect 149112 3408 149118 3460
rect 149514 3408 149520 3460
rect 149572 3448 149578 3460
rect 156046 3448 156052 3460
rect 149572 3420 156052 3448
rect 149572 3408 149578 3420
rect 156046 3408 156052 3420
rect 156104 3408 156110 3460
rect 161290 3408 161296 3460
rect 161348 3448 161354 3460
rect 167086 3448 167092 3460
rect 161348 3420 167092 3448
rect 161348 3408 161354 3420
rect 167086 3408 167092 3420
rect 167144 3408 167150 3460
rect 175458 3408 175464 3460
rect 175516 3448 175522 3460
rect 179414 3448 179420 3460
rect 175516 3420 179420 3448
rect 175516 3408 175522 3420
rect 179414 3408 179420 3420
rect 179472 3408 179478 3460
rect 181438 3408 181444 3460
rect 181496 3448 181502 3460
rect 184934 3448 184940 3460
rect 181496 3420 184940 3448
rect 181496 3408 181502 3420
rect 184934 3408 184940 3420
rect 184992 3408 184998 3460
rect 190822 3408 190828 3460
rect 190880 3448 190886 3460
rect 194778 3448 194784 3460
rect 190880 3420 194784 3448
rect 190880 3408 190886 3420
rect 194778 3408 194784 3420
rect 194836 3408 194842 3460
rect 301314 3408 301320 3460
rect 301372 3448 301378 3460
rect 303154 3448 303160 3460
rect 301372 3420 303160 3448
rect 301372 3408 301378 3420
rect 303154 3408 303160 3420
rect 303212 3408 303218 3460
rect 307754 3408 307760 3460
rect 307812 3448 307818 3460
rect 311434 3448 311440 3460
rect 307812 3420 311440 3448
rect 307812 3408 307818 3420
rect 311434 3408 311440 3420
rect 311492 3408 311498 3460
rect 311526 3408 311532 3460
rect 311584 3448 311590 3460
rect 313826 3448 313832 3460
rect 311584 3420 313832 3448
rect 311584 3408 311590 3420
rect 313826 3408 313832 3420
rect 313884 3408 313890 3460
rect 317506 3408 317512 3460
rect 317564 3448 317570 3460
rect 322106 3448 322112 3460
rect 317564 3420 322112 3448
rect 317564 3408 317570 3420
rect 322106 3408 322112 3420
rect 322164 3408 322170 3460
rect 325050 3408 325056 3460
rect 325108 3448 325114 3460
rect 329190 3448 329196 3460
rect 325108 3420 329196 3448
rect 325108 3408 325114 3420
rect 329190 3408 329196 3420
rect 329248 3408 329254 3460
rect 329650 3408 329656 3460
rect 329708 3448 329714 3460
rect 333882 3448 333888 3460
rect 329708 3420 333888 3448
rect 329708 3408 329714 3420
rect 333882 3408 333888 3420
rect 333940 3408 333946 3460
rect 343726 3408 343732 3460
rect 343784 3448 343790 3460
rect 349246 3448 349252 3460
rect 343784 3420 349252 3448
rect 343784 3408 343790 3420
rect 349246 3408 349252 3420
rect 349304 3408 349310 3460
rect 351086 3408 351092 3460
rect 351144 3448 351150 3460
rect 357526 3448 357532 3460
rect 351144 3420 357532 3448
rect 351144 3408 351150 3420
rect 357526 3408 357532 3420
rect 357584 3408 357590 3460
rect 365714 3408 365720 3460
rect 365772 3448 365778 3460
rect 372890 3448 372896 3460
rect 365772 3420 372896 3448
rect 365772 3408 365778 3420
rect 372890 3408 372896 3420
rect 372948 3408 372954 3460
rect 373350 3408 373356 3460
rect 373408 3448 373414 3460
rect 381170 3448 381176 3460
rect 373408 3420 381176 3448
rect 373408 3408 373414 3420
rect 381170 3408 381176 3420
rect 381228 3408 381234 3460
rect 381722 3408 381728 3460
rect 381780 3448 381786 3460
rect 389450 3448 389456 3460
rect 381780 3420 389456 3448
rect 381780 3408 381786 3420
rect 389450 3408 389456 3420
rect 389508 3408 389514 3460
rect 390186 3408 390192 3460
rect 390244 3448 390250 3460
rect 397730 3448 397736 3460
rect 390244 3420 397736 3448
rect 390244 3408 390250 3420
rect 397730 3408 397736 3420
rect 397788 3408 397794 3460
rect 398742 3408 398748 3460
rect 398800 3448 398806 3460
rect 407206 3448 407212 3460
rect 398800 3420 407212 3448
rect 398800 3408 398806 3420
rect 407206 3408 407212 3420
rect 407264 3408 407270 3460
rect 414014 3408 414020 3460
rect 414072 3448 414078 3460
rect 414072 3420 419212 3448
rect 414072 3408 414078 3420
rect 13538 3340 13544 3392
rect 13596 3380 13602 3392
rect 23290 3380 23296 3392
rect 13596 3352 23296 3380
rect 13596 3340 13602 3352
rect 23290 3340 23296 3352
rect 23348 3340 23354 3392
rect 27706 3340 27712 3392
rect 27764 3380 27770 3392
rect 34698 3380 34704 3392
rect 27764 3352 34704 3380
rect 27764 3340 27770 3352
rect 34698 3340 34704 3352
rect 34756 3340 34762 3392
rect 65518 3340 65524 3392
rect 65576 3380 65582 3392
rect 72418 3380 72424 3392
rect 65576 3352 72424 3380
rect 65576 3340 65582 3352
rect 72418 3340 72424 3352
rect 72476 3340 72482 3392
rect 96246 3340 96252 3392
rect 96304 3380 96310 3392
rect 102134 3380 102140 3392
rect 96304 3352 102140 3380
rect 96304 3340 96310 3352
rect 102134 3340 102140 3352
rect 102192 3340 102198 3392
rect 115198 3340 115204 3392
rect 115256 3380 115262 3392
rect 122742 3380 122748 3392
rect 115256 3352 122748 3380
rect 115256 3340 115262 3352
rect 122742 3340 122748 3352
rect 122800 3340 122806 3392
rect 301866 3340 301872 3392
rect 301924 3380 301930 3392
rect 304350 3380 304356 3392
rect 301924 3352 304356 3380
rect 301924 3340 301930 3352
rect 304350 3340 304356 3352
rect 304408 3340 304414 3392
rect 335354 3340 335360 3392
rect 335412 3380 335418 3392
rect 340966 3380 340972 3392
rect 335412 3352 340972 3380
rect 335412 3340 335418 3352
rect 340966 3340 340972 3352
rect 341024 3340 341030 3392
rect 345106 3340 345112 3392
rect 345164 3380 345170 3392
rect 351638 3380 351644 3392
rect 345164 3352 351644 3380
rect 345164 3340 345170 3352
rect 351638 3340 351644 3352
rect 351696 3340 351702 3392
rect 393314 3340 393320 3392
rect 393372 3380 393378 3392
rect 402514 3380 402520 3392
rect 393372 3352 402520 3380
rect 393372 3340 393378 3352
rect 402514 3340 402520 3352
rect 402572 3340 402578 3392
rect 404354 3340 404360 3392
rect 404412 3380 404418 3392
rect 414290 3380 414296 3392
rect 404412 3352 414296 3380
rect 404412 3340 404418 3352
rect 414290 3340 414296 3352
rect 414348 3340 414354 3392
rect 417970 3340 417976 3392
rect 418028 3380 418034 3392
rect 419184 3380 419212 3420
rect 419442 3408 419448 3460
rect 419500 3448 419506 3460
rect 429654 3448 429660 3460
rect 419500 3420 429660 3448
rect 419500 3408 419506 3420
rect 429654 3408 429660 3420
rect 429712 3408 429718 3460
rect 433334 3408 433340 3460
rect 433392 3448 433398 3460
rect 445018 3448 445024 3460
rect 433392 3420 445024 3448
rect 433392 3408 433398 3420
rect 445018 3408 445024 3420
rect 445076 3408 445082 3460
rect 481634 3408 481640 3460
rect 481692 3448 481698 3460
rect 484026 3448 484032 3460
rect 481692 3420 484032 3448
rect 481692 3408 481698 3420
rect 484026 3408 484032 3420
rect 484084 3408 484090 3460
rect 487154 3408 487160 3460
rect 487212 3448 487218 3460
rect 489914 3448 489920 3460
rect 487212 3420 489920 3448
rect 487212 3408 487218 3420
rect 489914 3408 489920 3420
rect 489972 3408 489978 3460
rect 501046 3408 501052 3460
rect 501104 3448 501110 3460
rect 505370 3448 505376 3460
rect 501104 3420 505376 3448
rect 501104 3408 501110 3420
rect 505370 3408 505376 3420
rect 505428 3408 505434 3460
rect 506474 3408 506480 3460
rect 506532 3448 506538 3460
rect 510062 3448 510068 3460
rect 506532 3420 510068 3448
rect 506532 3408 506538 3420
rect 510062 3408 510068 3420
rect 510120 3408 510126 3460
rect 510706 3408 510712 3460
rect 510764 3448 510770 3460
rect 514754 3448 514760 3460
rect 510764 3420 514760 3448
rect 510764 3408 510770 3420
rect 514754 3408 514760 3420
rect 514812 3408 514818 3460
rect 517606 3408 517612 3460
rect 517664 3448 517670 3460
rect 523034 3448 523040 3460
rect 517664 3420 523040 3448
rect 517664 3408 517670 3420
rect 523034 3408 523040 3420
rect 523092 3408 523098 3460
rect 532602 3408 532608 3460
rect 532660 3448 532666 3460
rect 537202 3448 537208 3460
rect 532660 3420 537208 3448
rect 532660 3408 532666 3420
rect 537202 3408 537208 3420
rect 537260 3408 537266 3460
rect 543706 3448 543734 3488
rect 551922 3476 551928 3528
rect 551980 3516 551986 3528
rect 557350 3516 557356 3528
rect 551980 3488 557356 3516
rect 551980 3476 551986 3488
rect 557350 3476 557356 3488
rect 557408 3476 557414 3528
rect 572714 3516 572720 3528
rect 557460 3488 572720 3516
rect 552658 3448 552664 3460
rect 543706 3420 552664 3448
rect 552658 3408 552664 3420
rect 552716 3408 552722 3460
rect 552750 3408 552756 3460
rect 552808 3448 552814 3460
rect 557460 3448 557488 3488
rect 572714 3476 572720 3488
rect 572772 3476 572778 3528
rect 552808 3420 557488 3448
rect 552808 3408 552814 3420
rect 557534 3408 557540 3460
rect 557592 3448 557598 3460
rect 579798 3448 579804 3460
rect 557592 3420 579804 3448
rect 557592 3408 557598 3420
rect 579798 3408 579804 3420
rect 579856 3408 579862 3460
rect 424962 3380 424968 3392
rect 418028 3352 419120 3380
rect 419184 3352 424968 3380
rect 418028 3340 418034 3352
rect 8754 3272 8760 3324
rect 8812 3312 8818 3324
rect 17954 3312 17960 3324
rect 8812 3284 17960 3312
rect 8812 3272 8818 3284
rect 17954 3272 17960 3284
rect 18012 3272 18018 3324
rect 20622 3272 20628 3324
rect 20680 3312 20686 3324
rect 26326 3312 26332 3324
rect 20680 3284 26332 3312
rect 20680 3272 20686 3284
rect 26326 3272 26332 3284
rect 26384 3272 26390 3324
rect 40678 3272 40684 3324
rect 40736 3312 40742 3324
rect 46934 3312 46940 3324
rect 40736 3284 46940 3312
rect 40736 3272 40742 3284
rect 46934 3272 46940 3284
rect 46992 3272 46998 3324
rect 48958 3272 48964 3324
rect 49016 3312 49022 3324
rect 55214 3312 55220 3324
rect 49016 3284 55220 3312
rect 49016 3272 49022 3284
rect 55214 3272 55220 3284
rect 55272 3272 55278 3324
rect 78582 3272 78588 3324
rect 78640 3312 78646 3324
rect 84286 3312 84292 3324
rect 78640 3284 84292 3312
rect 78640 3272 78646 3284
rect 84286 3272 84292 3284
rect 84344 3272 84350 3324
rect 87966 3272 87972 3324
rect 88024 3312 88030 3324
rect 93854 3312 93860 3324
rect 88024 3284 93860 3312
rect 88024 3272 88030 3284
rect 93854 3272 93860 3284
rect 93912 3272 93918 3324
rect 117590 3272 117596 3324
rect 117648 3312 117654 3324
rect 124214 3312 124220 3324
rect 117648 3284 124220 3312
rect 117648 3272 117654 3284
rect 124214 3272 124220 3284
rect 124272 3272 124278 3324
rect 143534 3272 143540 3324
rect 143592 3312 143598 3324
rect 150434 3312 150440 3324
rect 143592 3284 150440 3312
rect 143592 3272 143598 3284
rect 150434 3272 150440 3284
rect 150492 3272 150498 3324
rect 154206 3272 154212 3324
rect 154264 3312 154270 3324
rect 160186 3312 160192 3324
rect 154264 3284 160192 3312
rect 154264 3272 154270 3284
rect 160186 3272 160192 3284
rect 160244 3272 160250 3324
rect 162486 3272 162492 3324
rect 162544 3312 162550 3324
rect 166994 3312 167000 3324
rect 162544 3284 167000 3312
rect 162544 3272 162550 3284
rect 166994 3272 167000 3284
rect 167052 3272 167058 3324
rect 176654 3272 176660 3324
rect 176712 3312 176718 3324
rect 180794 3312 180800 3324
rect 176712 3284 180800 3312
rect 176712 3272 176718 3284
rect 180794 3272 180800 3284
rect 180852 3272 180858 3324
rect 186130 3272 186136 3324
rect 186188 3312 186194 3324
rect 189166 3312 189172 3324
rect 186188 3284 189172 3312
rect 186188 3272 186194 3284
rect 189166 3272 189172 3284
rect 189224 3272 189230 3324
rect 194410 3272 194416 3324
rect 194468 3312 194474 3324
rect 197446 3312 197452 3324
rect 194468 3284 197452 3312
rect 194468 3272 194474 3284
rect 197446 3272 197452 3284
rect 197504 3272 197510 3324
rect 202690 3272 202696 3324
rect 202748 3312 202754 3324
rect 205726 3312 205732 3324
rect 202748 3284 205732 3312
rect 202748 3272 202754 3284
rect 205726 3272 205732 3284
rect 205784 3272 205790 3324
rect 296714 3272 296720 3324
rect 296772 3312 296778 3324
rect 299658 3312 299664 3324
rect 296772 3284 299664 3312
rect 296772 3272 296778 3284
rect 299658 3272 299664 3284
rect 299716 3272 299722 3324
rect 306466 3272 306472 3324
rect 306524 3312 306530 3324
rect 310238 3312 310244 3324
rect 306524 3284 310244 3312
rect 306524 3272 306530 3284
rect 310238 3272 310244 3284
rect 310296 3272 310302 3324
rect 314562 3272 314568 3324
rect 314620 3312 314626 3324
rect 317322 3312 317328 3324
rect 314620 3284 317328 3312
rect 314620 3272 314626 3284
rect 317322 3272 317328 3284
rect 317380 3272 317386 3324
rect 317414 3272 317420 3324
rect 317472 3312 317478 3324
rect 320910 3312 320916 3324
rect 317472 3284 320916 3312
rect 317472 3272 317478 3284
rect 320910 3272 320916 3284
rect 320968 3272 320974 3324
rect 326246 3272 326252 3324
rect 326304 3312 326310 3324
rect 330386 3312 330392 3324
rect 326304 3284 330392 3312
rect 326304 3272 326310 3284
rect 330386 3272 330392 3284
rect 330444 3272 330450 3324
rect 331122 3272 331128 3324
rect 331180 3312 331186 3324
rect 335078 3312 335084 3324
rect 331180 3284 335084 3312
rect 331180 3272 331186 3284
rect 335078 3272 335084 3284
rect 335136 3272 335142 3324
rect 339402 3272 339408 3324
rect 339460 3312 339466 3324
rect 343358 3312 343364 3324
rect 339460 3284 343364 3312
rect 339460 3272 339466 3284
rect 343358 3272 343364 3284
rect 343416 3272 343422 3324
rect 345014 3272 345020 3324
rect 345072 3312 345078 3324
rect 350442 3312 350448 3324
rect 345072 3284 350448 3312
rect 345072 3272 345078 3284
rect 350442 3272 350448 3284
rect 350500 3272 350506 3324
rect 379330 3272 379336 3324
rect 379388 3312 379394 3324
rect 385954 3312 385960 3324
rect 379388 3284 385960 3312
rect 379388 3272 379394 3284
rect 385954 3272 385960 3284
rect 386012 3272 386018 3324
rect 408494 3272 408500 3324
rect 408552 3312 408558 3324
rect 418982 3312 418988 3324
rect 408552 3284 418988 3312
rect 408552 3272 408558 3284
rect 418982 3272 418988 3284
rect 419040 3272 419046 3324
rect 419092 3312 419120 3352
rect 424962 3340 424968 3352
rect 425020 3340 425026 3392
rect 513190 3340 513196 3392
rect 513248 3380 513254 3392
rect 517146 3380 517152 3392
rect 513248 3352 517152 3380
rect 513248 3340 513254 3352
rect 517146 3340 517152 3352
rect 517204 3340 517210 3392
rect 520458 3340 520464 3392
rect 520516 3380 520522 3392
rect 525426 3380 525432 3392
rect 520516 3352 525432 3380
rect 520516 3340 520522 3352
rect 525426 3340 525432 3352
rect 525484 3340 525490 3392
rect 530026 3340 530032 3392
rect 530084 3380 530090 3392
rect 536098 3380 536104 3392
rect 530084 3352 536104 3380
rect 530084 3340 530090 3352
rect 536098 3340 536104 3352
rect 536156 3340 536162 3392
rect 545114 3340 545120 3392
rect 545172 3380 545178 3392
rect 545172 3352 552704 3380
rect 545172 3340 545178 3352
rect 427262 3312 427268 3324
rect 419092 3284 427268 3312
rect 427262 3272 427268 3284
rect 427320 3272 427326 3324
rect 500954 3272 500960 3324
rect 501012 3312 501018 3324
rect 504174 3312 504180 3324
rect 501012 3284 504180 3312
rect 501012 3272 501018 3284
rect 504174 3272 504180 3284
rect 504232 3272 504238 3324
rect 510154 3272 510160 3324
rect 510212 3312 510218 3324
rect 513558 3312 513564 3324
rect 510212 3284 513564 3312
rect 510212 3272 510218 3284
rect 513558 3272 513564 3284
rect 513616 3272 513622 3324
rect 135254 3204 135260 3256
rect 135312 3244 135318 3256
rect 142154 3244 142160 3256
rect 135312 3216 142160 3244
rect 135312 3204 135318 3216
rect 142154 3204 142160 3216
rect 142212 3204 142218 3256
rect 164878 3204 164884 3256
rect 164936 3244 164942 3256
rect 169754 3244 169760 3256
rect 164936 3216 169760 3244
rect 164936 3204 164942 3216
rect 169754 3204 169760 3216
rect 169812 3204 169818 3256
rect 184934 3204 184940 3256
rect 184992 3244 184998 3256
rect 189074 3244 189080 3256
rect 184992 3216 189080 3244
rect 184992 3204 184998 3216
rect 189074 3204 189080 3216
rect 189132 3204 189138 3256
rect 195606 3204 195612 3256
rect 195664 3244 195670 3256
rect 198826 3244 198832 3256
rect 195664 3216 198832 3244
rect 195664 3204 195670 3216
rect 198826 3204 198832 3216
rect 198884 3204 198890 3256
rect 320082 3204 320088 3256
rect 320140 3244 320146 3256
rect 323302 3244 323308 3256
rect 320140 3216 323308 3244
rect 320140 3204 320146 3216
rect 323302 3204 323308 3216
rect 323360 3204 323366 3256
rect 340782 3204 340788 3256
rect 340840 3244 340846 3256
rect 344554 3244 344560 3256
rect 340840 3216 344560 3244
rect 340840 3204 340846 3216
rect 344554 3204 344560 3216
rect 344612 3204 344618 3256
rect 356054 3204 356060 3256
rect 356112 3244 356118 3256
rect 363506 3244 363512 3256
rect 356112 3216 363512 3244
rect 356112 3204 356118 3216
rect 363506 3204 363512 3216
rect 363564 3204 363570 3256
rect 503622 3204 503628 3256
rect 503680 3244 503686 3256
rect 506474 3244 506480 3256
rect 503680 3216 506480 3244
rect 503680 3204 503686 3216
rect 506474 3204 506480 3216
rect 506532 3204 506538 3256
rect 518894 3204 518900 3256
rect 518952 3244 518958 3256
rect 524230 3244 524236 3256
rect 518952 3216 524236 3244
rect 518952 3204 518958 3216
rect 524230 3204 524236 3216
rect 524288 3204 524294 3256
rect 540974 3204 540980 3256
rect 541032 3244 541038 3256
rect 547874 3244 547880 3256
rect 541032 3216 547880 3244
rect 541032 3204 541038 3216
rect 547874 3204 547880 3216
rect 547932 3204 547938 3256
rect 552676 3244 552704 3352
rect 557626 3340 557632 3392
rect 557684 3380 557690 3392
rect 565630 3380 565636 3392
rect 557684 3352 565636 3380
rect 557684 3340 557690 3352
rect 565630 3340 565636 3352
rect 565688 3340 565694 3392
rect 553210 3272 553216 3324
rect 553268 3312 553274 3324
rect 573910 3312 573916 3324
rect 553268 3284 573916 3312
rect 553268 3272 553274 3284
rect 573910 3272 573916 3284
rect 573968 3272 573974 3324
rect 566826 3244 566832 3256
rect 552676 3216 566832 3244
rect 566826 3204 566832 3216
rect 566884 3204 566890 3256
rect 17034 3136 17040 3188
rect 17092 3176 17098 3188
rect 24026 3176 24032 3188
rect 17092 3148 24032 3176
rect 17092 3136 17098 3148
rect 24026 3136 24032 3148
rect 24084 3136 24090 3188
rect 98638 3136 98644 3188
rect 98696 3176 98702 3188
rect 104986 3176 104992 3188
rect 98696 3148 104992 3176
rect 98696 3136 98702 3148
rect 104986 3136 104992 3148
rect 105044 3136 105050 3188
rect 126974 3136 126980 3188
rect 127032 3176 127038 3188
rect 133966 3176 133972 3188
rect 127032 3148 133972 3176
rect 127032 3136 127038 3148
rect 133966 3136 133972 3148
rect 134024 3136 134030 3188
rect 173158 3136 173164 3188
rect 173216 3176 173222 3188
rect 178034 3176 178040 3188
rect 173216 3148 178040 3176
rect 173216 3136 173222 3148
rect 178034 3136 178040 3148
rect 178092 3136 178098 3188
rect 182542 3136 182548 3188
rect 182600 3176 182606 3188
rect 186314 3176 186320 3188
rect 182600 3148 186320 3176
rect 182600 3136 182606 3148
rect 186314 3136 186320 3148
rect 186372 3136 186378 3188
rect 291654 3136 291660 3188
rect 291712 3176 291718 3188
rect 293678 3176 293684 3188
rect 291712 3148 293684 3176
rect 291712 3136 291718 3148
rect 293678 3136 293684 3148
rect 293736 3136 293742 3188
rect 298094 3136 298100 3188
rect 298152 3176 298158 3188
rect 300762 3176 300768 3188
rect 298152 3148 300768 3176
rect 298152 3136 298158 3148
rect 300762 3136 300768 3148
rect 300820 3136 300826 3188
rect 312722 3136 312728 3188
rect 312780 3176 312786 3188
rect 315022 3176 315028 3188
rect 312780 3148 315028 3176
rect 312780 3136 312786 3148
rect 315022 3136 315028 3148
rect 315080 3136 315086 3188
rect 321462 3136 321468 3188
rect 321520 3176 321526 3188
rect 324406 3176 324412 3188
rect 321520 3148 324412 3176
rect 321520 3136 321526 3148
rect 324406 3136 324412 3148
rect 324464 3136 324470 3188
rect 327074 3136 327080 3188
rect 327132 3176 327138 3188
rect 331582 3176 331588 3188
rect 327132 3148 331588 3176
rect 327132 3136 327138 3148
rect 331582 3136 331588 3148
rect 331640 3136 331646 3188
rect 486326 3136 486332 3188
rect 486384 3176 486390 3188
rect 488810 3176 488816 3188
rect 486384 3148 488816 3176
rect 486384 3136 486390 3148
rect 488810 3136 488816 3148
rect 488868 3136 488874 3188
rect 490006 3136 490012 3188
rect 490064 3176 490070 3188
rect 493502 3176 493508 3188
rect 490064 3148 493508 3176
rect 490064 3136 490070 3148
rect 493502 3136 493508 3148
rect 493560 3136 493566 3188
rect 495526 3136 495532 3188
rect 495584 3176 495590 3188
rect 498194 3176 498200 3188
rect 495584 3148 498200 3176
rect 495584 3136 495590 3148
rect 498194 3136 498200 3148
rect 498252 3136 498258 3188
rect 505002 3136 505008 3188
rect 505060 3176 505066 3188
rect 507670 3176 507676 3188
rect 505060 3148 507676 3176
rect 505060 3136 505066 3148
rect 507670 3136 507676 3148
rect 507728 3136 507734 3188
rect 514662 3136 514668 3188
rect 514720 3176 514726 3188
rect 518342 3176 518348 3188
rect 514720 3148 518348 3176
rect 514720 3136 514726 3148
rect 518342 3136 518348 3148
rect 518400 3136 518406 3188
rect 522942 3136 522948 3188
rect 523000 3176 523006 3188
rect 526622 3176 526628 3188
rect 523000 3148 526628 3176
rect 523000 3136 523006 3148
rect 526622 3136 526628 3148
rect 526680 3136 526686 3188
rect 555418 3136 555424 3188
rect 555476 3176 555482 3188
rect 562042 3176 562048 3188
rect 555476 3148 562048 3176
rect 555476 3136 555482 3148
rect 562042 3136 562048 3148
rect 562100 3136 562106 3188
rect 374362 3068 374368 3120
rect 374420 3108 374426 3120
rect 382366 3108 382372 3120
rect 374420 3080 382372 3108
rect 374420 3068 374426 3080
rect 382366 3068 382372 3080
rect 382424 3068 382430 3120
rect 38378 3000 38384 3052
rect 38436 3040 38442 3052
rect 44358 3040 44364 3052
rect 38436 3012 44364 3040
rect 38436 3000 38442 3012
rect 44358 3000 44364 3012
rect 44416 3000 44422 3052
rect 76190 3000 76196 3052
rect 76248 3040 76254 3052
rect 82814 3040 82820 3052
rect 76248 3012 82820 3040
rect 76248 3000 76254 3012
rect 82814 3000 82820 3012
rect 82872 3000 82878 3052
rect 84470 3000 84476 3052
rect 84528 3040 84534 3052
rect 91186 3040 91192 3052
rect 84528 3012 91192 3040
rect 84528 3000 84534 3012
rect 91186 3000 91192 3012
rect 91244 3000 91250 3052
rect 114002 3000 114008 3052
rect 114060 3040 114066 3052
rect 120166 3040 120172 3052
rect 114060 3012 120172 3040
rect 114060 3000 114066 3012
rect 120166 3000 120172 3012
rect 120224 3000 120230 3052
rect 123478 3000 123484 3052
rect 123536 3040 123542 3052
rect 131022 3040 131028 3052
rect 123536 3012 131028 3040
rect 123536 3000 123542 3012
rect 131022 3000 131028 3012
rect 131080 3000 131086 3052
rect 134150 3000 134156 3052
rect 134208 3040 134214 3052
rect 140774 3040 140780 3052
rect 134208 3012 140780 3040
rect 134208 3000 134214 3012
rect 140774 3000 140780 3012
rect 140832 3000 140838 3052
rect 144730 3000 144736 3052
rect 144788 3040 144794 3052
rect 150526 3040 150532 3052
rect 144788 3012 150532 3040
rect 144788 3000 144794 3012
rect 150526 3000 150532 3012
rect 150584 3000 150590 3052
rect 278774 3000 278780 3052
rect 278832 3040 278838 3052
rect 280706 3040 280712 3052
rect 278832 3012 280712 3040
rect 278832 3000 278838 3012
rect 280706 3000 280712 3012
rect 280764 3000 280770 3052
rect 284662 3000 284668 3052
rect 284720 3040 284726 3052
rect 286594 3040 286600 3052
rect 284720 3012 286600 3040
rect 284720 3000 284726 3012
rect 286594 3000 286600 3012
rect 286652 3000 286658 3052
rect 288434 3000 288440 3052
rect 288492 3040 288498 3052
rect 290182 3040 290188 3052
rect 288492 3012 290188 3040
rect 288492 3000 288498 3012
rect 290182 3000 290188 3012
rect 290240 3000 290246 3052
rect 294230 3000 294236 3052
rect 294288 3040 294294 3052
rect 296070 3040 296076 3052
rect 294288 3012 296076 3040
rect 294288 3000 294294 3012
rect 296070 3000 296076 3012
rect 296128 3000 296134 3052
rect 356146 3000 356152 3052
rect 356204 3040 356210 3052
rect 362310 3040 362316 3052
rect 356204 3012 362316 3040
rect 356204 3000 356210 3012
rect 362310 3000 362316 3012
rect 362368 3000 362374 3052
rect 364794 3000 364800 3052
rect 364852 3040 364858 3052
rect 371694 3040 371700 3052
rect 364852 3012 371700 3040
rect 364852 3000 364858 3012
rect 371694 3000 371700 3012
rect 371752 3000 371758 3052
rect 383654 3000 383660 3052
rect 383712 3040 383718 3052
rect 393038 3040 393044 3052
rect 383712 3012 393044 3040
rect 383712 3000 383718 3012
rect 393038 3000 393044 3012
rect 393096 3000 393102 3052
rect 475102 3000 475108 3052
rect 475160 3040 475166 3052
rect 476942 3040 476948 3052
rect 475160 3012 476948 3040
rect 475160 3000 475166 3012
rect 476942 3000 476948 3012
rect 477000 3000 477006 3052
rect 485682 3000 485688 3052
rect 485740 3040 485746 3052
rect 487614 3040 487620 3052
rect 485740 3012 487620 3040
rect 485740 3000 485746 3012
rect 487614 3000 487620 3012
rect 487672 3000 487678 3052
rect 493962 3000 493968 3052
rect 494020 3040 494026 3052
rect 495894 3040 495900 3052
rect 494020 3012 495900 3040
rect 494020 3000 494026 3012
rect 495894 3000 495900 3012
rect 495952 3000 495958 3052
rect 496906 3000 496912 3052
rect 496964 3040 496970 3052
rect 500586 3040 500592 3052
rect 496964 3012 500592 3040
rect 496964 3000 496970 3012
rect 500586 3000 500592 3012
rect 500644 3000 500650 3052
rect 28902 2932 28908 2984
rect 28960 2972 28966 2984
rect 34882 2972 34888 2984
rect 28960 2944 34888 2972
rect 28960 2932 28966 2944
rect 34882 2932 34888 2944
rect 34940 2932 34946 2984
rect 35986 2932 35992 2984
rect 36044 2972 36050 2984
rect 43346 2972 43352 2984
rect 36044 2944 43352 2972
rect 36044 2932 36050 2944
rect 43346 2932 43352 2944
rect 43404 2932 43410 2984
rect 46658 2932 46664 2984
rect 46716 2972 46722 2984
rect 53098 2972 53104 2984
rect 46716 2944 53104 2972
rect 46716 2932 46722 2944
rect 53098 2932 53104 2944
rect 53156 2932 53162 2984
rect 56042 2932 56048 2984
rect 56100 2972 56106 2984
rect 62666 2972 62672 2984
rect 56100 2944 62672 2972
rect 56100 2932 56106 2944
rect 62666 2932 62672 2944
rect 62724 2932 62730 2984
rect 66714 2932 66720 2984
rect 66772 2972 66778 2984
rect 73154 2972 73160 2984
rect 66772 2944 73160 2972
rect 66772 2932 66778 2944
rect 73154 2932 73160 2944
rect 73212 2932 73218 2984
rect 124674 2932 124680 2984
rect 124732 2972 124738 2984
rect 132402 2972 132408 2984
rect 124732 2944 132408 2972
rect 124732 2932 124738 2944
rect 132402 2932 132408 2944
rect 132460 2932 132466 2984
rect 132954 2932 132960 2984
rect 133012 2972 133018 2984
rect 139578 2972 139584 2984
rect 133012 2944 139584 2972
rect 133012 2932 133018 2944
rect 139578 2932 139584 2944
rect 139636 2932 139642 2984
rect 147122 2932 147128 2984
rect 147180 2972 147186 2984
rect 153194 2972 153200 2984
rect 147180 2944 153200 2972
rect 147180 2932 147186 2944
rect 153194 2932 153200 2944
rect 153252 2932 153258 2984
rect 156598 2932 156604 2984
rect 156656 2972 156662 2984
rect 161474 2972 161480 2984
rect 156656 2944 161480 2972
rect 156656 2932 156662 2944
rect 161474 2932 161480 2944
rect 161532 2932 161538 2984
rect 287238 2932 287244 2984
rect 287296 2972 287302 2984
rect 288986 2972 288992 2984
rect 287296 2944 288992 2972
rect 287296 2932 287302 2944
rect 288986 2932 288992 2944
rect 289044 2932 289050 2984
rect 375374 2932 375380 2984
rect 375432 2972 375438 2984
rect 383562 2972 383568 2984
rect 375432 2944 383568 2972
rect 375432 2932 375438 2944
rect 383562 2932 383568 2944
rect 383620 2932 383626 2984
rect 384390 2932 384396 2984
rect 384448 2972 384454 2984
rect 391842 2972 391848 2984
rect 384448 2944 391848 2972
rect 384448 2932 384454 2944
rect 391842 2932 391848 2944
rect 391900 2932 391906 2984
rect 484670 2932 484676 2984
rect 484728 2972 484734 2984
rect 486418 2972 486424 2984
rect 484728 2944 486424 2972
rect 484728 2932 484734 2944
rect 486418 2932 486424 2944
rect 486476 2932 486482 2984
rect 539686 2932 539692 2984
rect 539744 2972 539750 2984
rect 545482 2972 545488 2984
rect 539744 2944 545488 2972
rect 539744 2932 539750 2944
rect 545482 2932 545488 2944
rect 545540 2932 545546 2984
rect 86862 2864 86868 2916
rect 86920 2904 86926 2916
rect 92474 2904 92480 2916
rect 86920 2876 92480 2904
rect 86920 2864 86926 2876
rect 92474 2864 92480 2876
rect 92532 2864 92538 2916
rect 93946 2864 93952 2916
rect 94004 2904 94010 2916
rect 100938 2904 100944 2916
rect 94004 2876 100944 2904
rect 94004 2864 94010 2876
rect 100938 2864 100944 2876
rect 100996 2864 101002 2916
rect 105722 2864 105728 2916
rect 105780 2904 105786 2916
rect 111978 2904 111984 2916
rect 105780 2876 111984 2904
rect 105780 2864 105786 2876
rect 111978 2864 111984 2876
rect 112036 2864 112042 2916
rect 153010 2864 153016 2916
rect 153068 2904 153074 2916
rect 158714 2904 158720 2916
rect 153068 2876 158720 2904
rect 153068 2864 153074 2876
rect 158714 2864 158720 2876
rect 158772 2864 158778 2916
rect 336734 2864 336740 2916
rect 336792 2904 336798 2916
rect 342162 2904 342168 2916
rect 336792 2876 342168 2904
rect 336792 2864 336798 2876
rect 342162 2864 342168 2876
rect 342220 2864 342226 2916
rect 349062 2864 349068 2916
rect 349120 2904 349126 2916
rect 354030 2904 354036 2916
rect 349120 2876 354036 2904
rect 349120 2864 349126 2876
rect 354030 2864 354036 2876
rect 354088 2864 354094 2916
rect 495342 2864 495348 2916
rect 495400 2904 495406 2916
rect 497090 2904 497096 2916
rect 495400 2876 497096 2904
rect 495400 2864 495406 2876
rect 497090 2864 497096 2876
rect 497148 2864 497154 2916
rect 528646 2864 528652 2916
rect 528704 2904 528710 2916
rect 534902 2904 534908 2916
rect 528704 2876 534908 2904
rect 528704 2864 528710 2876
rect 534902 2864 534908 2876
rect 534960 2864 534966 2916
<< via1 >>
rect 71780 702992 71832 703044
rect 72976 702992 73028 703044
rect 527272 700476 527324 700528
rect 543464 700476 543516 700528
rect 495440 700408 495492 700460
rect 510988 700408 511040 700460
rect 542360 700340 542412 700392
rect 559656 700340 559708 700392
rect 342260 700272 342312 700324
rect 348792 700272 348844 700324
rect 372620 700272 372672 700324
rect 381176 700272 381228 700324
rect 387800 700272 387852 700324
rect 397460 700272 397512 700324
rect 402980 700272 403032 700324
rect 413652 700272 413704 700324
rect 419540 700272 419592 700324
rect 429844 700272 429896 700324
rect 434720 700272 434772 700324
rect 446128 700272 446180 700324
rect 449900 700272 449952 700324
rect 462320 700272 462372 700324
rect 465080 700272 465132 700324
rect 478512 700272 478564 700324
rect 480260 700272 480312 700324
rect 494796 700272 494848 700324
rect 510620 700272 510672 700324
rect 527180 700272 527232 700324
rect 557540 700272 557592 700324
rect 575848 700272 575900 700324
rect 105452 699728 105504 699780
rect 108304 699728 108356 699780
rect 121644 699660 121696 699712
rect 124864 699660 124916 699712
rect 137836 699660 137888 699712
rect 140044 699660 140096 699712
rect 154120 699660 154172 699712
rect 156604 699660 156656 699712
rect 170312 699660 170364 699712
rect 172520 699660 172572 699712
rect 186504 699660 186556 699712
rect 189080 699660 189132 699712
rect 202788 699660 202840 699712
rect 204260 699660 204312 699712
rect 249800 699660 249852 699712
rect 251456 699660 251508 699712
rect 264980 699660 265032 699712
rect 267648 699660 267700 699712
rect 280160 699660 280212 699712
rect 283840 699660 283892 699712
rect 296720 699660 296772 699712
rect 300124 699660 300176 699712
rect 311900 699660 311952 699712
rect 316316 699660 316368 699712
rect 327080 699660 327132 699712
rect 332508 699660 332560 699712
rect 569224 696940 569276 696992
rect 580172 696940 580224 696992
rect 569316 683136 569368 683188
rect 580172 683136 580224 683188
rect 6920 680960 6972 681012
rect 19892 680960 19944 681012
rect 23480 680960 23532 681012
rect 35256 680960 35308 681012
rect 40040 680960 40092 681012
rect 50620 680960 50672 681012
rect 56600 680960 56652 681012
rect 66260 680960 66312 681012
rect 71780 680960 71832 681012
rect 81440 680960 81492 681012
rect 88340 680960 88392 681012
rect 96712 680960 96764 681012
rect 140044 680756 140096 680808
rect 142804 680756 142856 680808
rect 358544 680688 358596 680740
rect 364340 680688 364392 680740
rect 108304 680552 108356 680604
rect 112076 680552 112128 680604
rect 156604 680552 156656 680604
rect 158168 680552 158220 680604
rect 218060 680552 218112 680604
rect 219716 680552 219768 680604
rect 124864 680416 124916 680468
rect 127440 680416 127492 680468
rect 569408 670692 569460 670744
rect 580172 670692 580224 670744
rect 3424 670624 3476 670676
rect 9404 670624 9456 670676
rect 3516 658180 3568 658232
rect 9404 658180 9456 658232
rect 569224 656888 569276 656940
rect 580172 656888 580224 656940
rect 3608 645804 3660 645856
rect 9404 645804 9456 645856
rect 569316 643084 569368 643136
rect 580172 643084 580224 643136
rect 3424 633360 3476 633412
rect 8668 633360 8720 633412
rect 569224 630640 569276 630692
rect 580172 630640 580224 630692
rect 3516 620916 3568 620968
rect 8668 620916 8720 620968
rect 569316 616836 569368 616888
rect 580172 616836 580224 616888
rect 3608 607928 3660 607980
rect 9404 607928 9456 607980
rect 569408 603100 569460 603152
rect 580172 603100 580224 603152
rect 3424 596096 3476 596148
rect 9404 596096 9456 596148
rect 2780 592016 2832 592068
rect 6276 592016 6328 592068
rect 569224 590656 569276 590708
rect 579804 590656 579856 590708
rect 3516 585080 3568 585132
rect 9404 585080 9456 585132
rect 2964 579640 3016 579692
rect 6184 579640 6236 579692
rect 569316 576852 569368 576904
rect 580172 576852 580224 576904
rect 6276 572636 6328 572688
rect 8852 572636 8904 572688
rect 569224 563048 569276 563100
rect 579804 563048 579856 563100
rect 6184 559784 6236 559836
rect 9404 559784 9456 559836
rect 569316 550604 569368 550656
rect 580172 550604 580224 550656
rect 3424 547816 3476 547868
rect 9404 547816 9456 547868
rect 3424 539588 3476 539640
rect 7656 539588 7708 539640
rect 569224 536800 569276 536852
rect 580172 536800 580224 536852
rect 3516 535372 3568 535424
rect 9404 535372 9456 535424
rect 3424 527144 3476 527196
rect 7564 527144 7616 527196
rect 569316 524424 569368 524476
rect 580172 524424 580224 524476
rect 3424 514768 3476 514820
rect 8944 514768 8996 514820
rect 569224 510620 569276 510672
rect 580172 510620 580224 510672
rect 3056 500964 3108 501016
rect 9036 500964 9088 501016
rect 577504 496816 577556 496868
rect 579896 496816 579948 496868
rect 3424 488656 3476 488708
rect 8944 488656 8996 488708
rect 577596 484372 577648 484424
rect 580632 484372 580684 484424
rect 569868 482944 569920 482996
rect 577504 482944 577556 482996
rect 3424 475600 3476 475652
rect 9036 475600 9088 475652
rect 576124 470568 576176 470620
rect 579988 470568 580040 470620
rect 569868 470500 569920 470552
rect 577596 470500 577648 470552
rect 3424 462544 3476 462596
rect 8944 462544 8996 462596
rect 569868 457852 569920 457904
rect 576124 457852 576176 457904
rect 2780 449420 2832 449472
rect 6276 449420 6328 449472
rect 569132 445680 569184 445732
rect 580264 445680 580316 445732
rect 6276 437384 6328 437436
rect 9404 437384 9456 437436
rect 2964 436160 3016 436212
rect 6184 436160 6236 436212
rect 569316 433236 569368 433288
rect 580356 433236 580408 433288
rect 569224 430584 569276 430636
rect 580172 430584 580224 430636
rect 6184 424396 6236 424448
rect 9404 424396 9456 424448
rect 3424 423172 3476 423224
rect 7564 423172 7616 423224
rect 569224 418140 569276 418192
rect 580172 418140 580224 418192
rect 3148 409844 3200 409896
rect 7564 409844 7616 409896
rect 574744 404336 574796 404388
rect 580172 404336 580224 404388
rect 3424 397468 3476 397520
rect 7564 397468 7616 397520
rect 569132 395768 569184 395820
rect 574744 395768 574796 395820
rect 3424 383800 3476 383852
rect 7564 383800 7616 383852
rect 569868 383596 569920 383648
rect 578884 383596 578936 383648
rect 3424 371288 3476 371340
rect 7564 371288 7616 371340
rect 569592 371152 569644 371204
rect 578884 371152 578936 371204
rect 578240 364692 578292 364744
rect 579620 364692 579672 364744
rect 569684 358708 569736 358760
rect 578240 358708 578292 358760
rect 2780 357688 2832 357740
rect 4804 357688 4856 357740
rect 4804 351840 4856 351892
rect 8668 351840 8720 351892
rect 569684 346332 569736 346384
rect 579528 346332 579580 346384
rect 4160 339396 4212 339448
rect 9404 339396 9456 339448
rect 569224 338104 569276 338156
rect 580172 338104 580224 338156
rect 3056 327020 3108 327072
rect 9404 327020 9456 327072
rect 568672 321512 568724 321564
rect 580172 321512 580224 321564
rect 3424 314576 3476 314628
rect 9404 314576 9456 314628
rect 568948 311856 569000 311908
rect 580172 311856 580224 311908
rect 3424 306144 3476 306196
rect 9404 306144 9456 306196
rect 569868 295264 569920 295316
rect 580356 295264 580408 295316
rect 3424 292544 3476 292596
rect 9404 292544 9456 292596
rect 572720 284316 572772 284368
rect 580172 284316 580224 284368
rect 569868 282684 569920 282736
rect 572720 282684 572772 282736
rect 3424 279692 3476 279744
rect 9220 279692 9272 279744
rect 572720 271872 572772 271924
rect 579804 271872 579856 271924
rect 569316 270172 569368 270224
rect 572720 270172 572772 270224
rect 3056 266364 3108 266416
rect 9404 266364 9456 266416
rect 569132 258000 569184 258052
rect 579712 258068 579764 258120
rect 3424 254056 3476 254108
rect 9404 254056 9456 254108
rect 568672 244876 568724 244928
rect 580172 244876 580224 244928
rect 3424 240864 3476 240916
rect 9404 240864 9456 240916
rect 569868 232500 569920 232552
rect 580172 232500 580224 232552
rect 3424 227944 3476 227996
rect 8852 227944 8904 227996
rect 569500 219444 569552 219496
rect 580448 219376 580500 219428
rect 3424 214956 3476 215008
rect 8208 214956 8260 215008
rect 569868 207000 569920 207052
rect 579528 207000 579580 207052
rect 3332 202172 3384 202224
rect 8208 202172 8260 202224
rect 569316 194556 569368 194608
rect 579528 194556 579580 194608
rect 3424 188844 3476 188896
rect 8208 188844 8260 188896
rect 569408 182180 569460 182232
rect 576860 182180 576912 182232
rect 576860 179324 576912 179376
rect 580264 179324 580316 179376
rect 3424 176604 3476 176656
rect 8208 176604 8260 176656
rect 569868 169736 569920 169788
rect 577964 169736 578016 169788
rect 577964 166948 578016 167000
rect 579988 166948 580040 167000
rect 3516 163344 3568 163396
rect 8208 163344 8260 163396
rect 569868 157360 569920 157412
rect 579528 157360 579580 157412
rect 3424 150356 3476 150408
rect 8944 150356 8996 150408
rect 569868 144916 569920 144968
rect 578884 144916 578936 144968
rect 3240 137912 3292 137964
rect 8300 137912 8352 137964
rect 569868 132472 569920 132524
rect 578240 132472 578292 132524
rect 4160 129752 4212 129804
rect 9036 129752 9088 129804
rect 578240 126896 578292 126948
rect 579620 126896 579672 126948
rect 4804 118668 4856 118720
rect 9404 118668 9456 118720
rect 568672 118668 568724 118720
rect 578884 118668 578936 118720
rect 2780 110712 2832 110764
rect 4804 110712 4856 110764
rect 4804 106292 4856 106344
rect 9404 106292 9456 106344
rect 569684 106292 569736 106344
rect 578884 106292 578936 106344
rect 2780 97724 2832 97776
rect 4804 97724 4856 97776
rect 569684 94392 569736 94444
rect 576124 94392 576176 94444
rect 4804 93848 4856 93900
rect 9404 93848 9456 93900
rect 576124 86912 576176 86964
rect 580172 86912 580224 86964
rect 2780 85212 2832 85264
rect 4804 85212 4856 85264
rect 569684 81404 569736 81456
rect 578884 81404 578936 81456
rect 3424 71612 3476 71664
rect 8944 71612 8996 71664
rect 569592 69028 569644 69080
rect 578884 69028 578936 69080
rect 3148 59168 3200 59220
rect 8944 59168 8996 59220
rect 4804 56584 4856 56636
rect 8852 56584 8904 56636
rect 569132 56584 569184 56636
rect 574744 56584 574796 56636
rect 574744 46860 574796 46912
rect 580172 46860 580224 46912
rect 2780 45500 2832 45552
rect 4804 45500 4856 45552
rect 4896 44140 4948 44192
rect 9404 44140 9456 44192
rect 569868 44140 569920 44192
rect 578884 44140 578936 44192
rect 2780 32852 2832 32904
rect 4896 32852 4948 32904
rect 4804 31764 4856 31816
rect 9036 31764 9088 31816
rect 569500 31764 569552 31816
rect 578976 31764 579028 31816
rect 2780 20340 2832 20392
rect 4804 20340 4856 20392
rect 569868 19320 569920 19372
rect 578884 19320 578936 19372
rect 75920 9596 75972 9648
rect 81716 9596 81768 9648
rect 122840 9596 122892 9648
rect 123668 9596 123720 9648
rect 229100 9596 229152 9648
rect 229652 9596 229704 9648
rect 448888 9596 448940 9648
rect 462780 9596 462832 9648
rect 463240 9596 463292 9648
rect 476304 9596 476356 9648
rect 478696 9596 478748 9648
rect 491392 9596 491444 9648
rect 501880 9596 501932 9648
rect 515956 9596 516008 9648
rect 518440 9596 518492 9648
rect 532608 9596 532660 9648
rect 26332 9528 26384 9580
rect 35348 9528 35400 9580
rect 35992 9528 36044 9580
rect 44180 9528 44232 9580
rect 68652 9528 68704 9580
rect 73988 9528 74040 9580
rect 78588 9528 78640 9580
rect 82820 9528 82872 9580
rect 103612 9528 103664 9580
rect 107108 9528 107160 9580
rect 109132 9528 109184 9580
rect 112628 9528 112680 9580
rect 124220 9528 124272 9580
rect 125876 9528 125928 9580
rect 203892 9528 203944 9580
rect 206468 9528 206520 9580
rect 271144 9528 271196 9580
rect 272432 9528 272484 9580
rect 321928 9528 321980 9580
rect 324228 9528 324280 9580
rect 338488 9528 338540 9580
rect 340788 9528 340840 9580
rect 381544 9528 381596 9580
rect 382924 9528 382976 9580
rect 410248 9528 410300 9580
rect 412364 9528 412416 9580
rect 445576 9528 445628 9580
rect 459192 9528 459244 9580
rect 467656 9528 467708 9580
rect 480628 9528 480680 9580
rect 482928 9528 482980 9580
rect 496452 9528 496504 9580
rect 499488 9528 499540 9580
rect 513196 9528 513248 9580
rect 516048 9528 516100 9580
rect 528652 9528 528704 9580
rect 535000 9528 535052 9580
rect 547880 9528 547932 9580
rect 17960 9460 18012 9512
rect 24308 9460 24360 9512
rect 26424 9460 26476 9512
rect 34520 9460 34572 9512
rect 34704 9460 34756 9512
rect 41972 9460 42024 9512
rect 45744 9460 45796 9512
rect 53012 9460 53064 9512
rect 68928 9460 68980 9512
rect 73160 9460 73212 9512
rect 76104 9460 76156 9512
rect 80612 9460 80664 9512
rect 84384 9460 84436 9512
rect 88340 9460 88392 9512
rect 93860 9460 93912 9512
rect 98276 9460 98328 9512
rect 98460 9460 98512 9512
rect 101588 9460 101640 9512
rect 104992 9460 105044 9512
rect 108212 9460 108264 9512
rect 109224 9460 109276 9512
rect 111800 9460 111852 9512
rect 114560 9460 114612 9512
rect 117320 9460 117372 9512
rect 118608 9460 118660 9512
rect 119252 9460 119304 9512
rect 124128 9460 124180 9512
rect 124772 9460 124824 9512
rect 129648 9460 129700 9512
rect 130292 9460 130344 9512
rect 155960 9460 156012 9512
rect 156788 9460 156840 9512
rect 161480 9460 161532 9512
rect 162308 9460 162360 9512
rect 167000 9460 167052 9512
rect 167828 9460 167880 9512
rect 172520 9460 172572 9512
rect 173348 9460 173400 9512
rect 192024 9460 192076 9512
rect 195428 9460 195480 9512
rect 200304 9460 200356 9512
rect 203156 9460 203208 9512
rect 206192 9460 206244 9512
rect 208676 9460 208728 9512
rect 209780 9460 209832 9512
rect 211988 9460 212040 9512
rect 214472 9460 214524 9512
rect 216680 9460 216732 9512
rect 216864 9460 216916 9512
rect 218612 9460 218664 9512
rect 220452 9460 220504 9512
rect 222200 9460 222252 9512
rect 222752 9460 222804 9512
rect 224132 9460 224184 9512
rect 226340 9460 226392 9512
rect 227720 9460 227772 9512
rect 235816 9460 235868 9512
rect 236276 9460 236328 9512
rect 256608 9460 256660 9512
rect 257068 9460 257120 9512
rect 259000 9460 259052 9512
rect 259552 9460 259604 9512
rect 262128 9460 262180 9512
rect 262956 9460 263008 9512
rect 264520 9460 264572 9512
rect 265348 9460 265400 9512
rect 270040 9460 270092 9512
rect 271236 9460 271288 9512
rect 273168 9460 273220 9512
rect 274548 9460 274600 9512
rect 277768 9460 277820 9512
rect 279516 9460 279568 9512
rect 279976 9460 280028 9512
rect 281448 9460 281500 9512
rect 284208 9460 284260 9512
rect 284668 9460 284720 9512
rect 287704 9460 287756 9512
rect 288440 9460 288492 9512
rect 290924 9460 290976 9512
rect 291660 9460 291712 9512
rect 293224 9460 293276 9512
rect 294236 9460 294288 9512
rect 295248 9460 295300 9512
rect 296260 9460 296312 9512
rect 297640 9460 297692 9512
rect 298100 9460 298152 9512
rect 299848 9460 299900 9512
rect 301320 9460 301372 9512
rect 303068 9460 303120 9512
rect 304448 9460 304500 9512
rect 308680 9460 308732 9512
rect 310428 9460 310480 9512
rect 311808 9460 311860 9512
rect 313188 9460 313240 9512
rect 314200 9460 314252 9512
rect 315856 9460 315908 9512
rect 319720 9460 319772 9512
rect 321468 9460 321520 9512
rect 322848 9460 322900 9512
rect 324136 9460 324188 9512
rect 325240 9460 325292 9512
rect 326252 9460 326304 9512
rect 327448 9460 327500 9512
rect 329748 9460 329800 9512
rect 330760 9460 330812 9512
rect 332508 9460 332560 9512
rect 336280 9460 336332 9512
rect 336740 9460 336792 9512
rect 339408 9460 339460 9512
rect 340696 9460 340748 9512
rect 341800 9460 341852 9512
rect 343548 9460 343600 9512
rect 347320 9460 347372 9512
rect 349068 9460 349120 9512
rect 350448 9460 350500 9512
rect 351092 9460 351144 9512
rect 351736 9460 351788 9512
rect 353208 9460 353260 9512
rect 355048 9460 355100 9512
rect 356152 9460 356204 9512
rect 357256 9460 357308 9512
rect 358728 9460 358780 9512
rect 366088 9460 366140 9512
rect 368388 9460 368440 9512
rect 370504 9460 370556 9512
rect 372160 9460 372212 9512
rect 372528 9460 372580 9512
rect 373356 9460 373408 9512
rect 376024 9460 376076 9512
rect 378048 9460 378100 9512
rect 380440 9460 380492 9512
rect 381728 9460 381780 9512
rect 385960 9460 386012 9512
rect 387708 9460 387760 9512
rect 389088 9460 389140 9512
rect 390468 9460 390520 9512
rect 391480 9460 391532 9512
rect 392492 9460 392544 9512
rect 397000 9460 397052 9512
rect 398748 9460 398800 9512
rect 400128 9460 400180 9512
rect 401416 9460 401468 9512
rect 406936 9460 406988 9512
rect 407396 9460 407448 9512
rect 408040 9460 408092 9512
rect 408500 9460 408552 9512
rect 409144 9460 409196 9512
rect 411168 9460 411220 9512
rect 413560 9460 413612 9512
rect 414020 9460 414072 9512
rect 416504 9460 416556 9512
rect 418068 9460 418120 9512
rect 419080 9460 419132 9512
rect 420828 9460 420880 9512
rect 426808 9460 426860 9512
rect 427820 9460 427872 9512
rect 444288 9460 444340 9512
rect 458088 9460 458140 9512
rect 469864 9460 469916 9512
rect 484308 9460 484360 9512
rect 486424 9460 486476 9512
rect 499672 9460 499724 9512
rect 502984 9460 503036 9512
rect 516508 9460 516560 9512
rect 528284 9460 528336 9512
rect 540980 9460 541032 9512
rect 24952 9392 25004 9444
rect 29828 9392 29880 9444
rect 33784 9392 33836 9444
rect 40868 9392 40920 9444
rect 41328 9392 41380 9444
rect 47492 9392 47544 9444
rect 52276 9392 52328 9444
rect 58532 9392 58584 9444
rect 59268 9392 59320 9444
rect 64052 9392 64104 9444
rect 66352 9392 66404 9444
rect 71780 9392 71832 9444
rect 74632 9392 74684 9444
rect 79508 9392 79560 9444
rect 89628 9392 89680 9444
rect 92756 9392 92808 9444
rect 99472 9392 99524 9444
rect 102692 9392 102744 9444
rect 106832 9392 106884 9444
rect 109316 9392 109368 9444
rect 113272 9392 113324 9444
rect 115940 9392 115992 9444
rect 117228 9392 117280 9444
rect 118148 9392 118200 9444
rect 118700 9392 118752 9444
rect 121460 9392 121512 9444
rect 128268 9392 128320 9444
rect 129188 9392 129240 9444
rect 193220 9392 193272 9444
rect 196532 9392 196584 9444
rect 205088 9392 205140 9444
rect 207572 9392 207624 9444
rect 213368 9392 213420 9444
rect 215300 9392 215352 9444
rect 215668 9392 215720 9444
rect 217508 9392 217560 9444
rect 221556 9392 221608 9444
rect 223028 9392 223080 9444
rect 225144 9392 225196 9444
rect 226432 9392 226484 9444
rect 227536 9392 227588 9444
rect 228548 9392 228600 9444
rect 272248 9392 272300 9444
rect 273628 9392 273680 9444
rect 274456 9392 274508 9444
rect 275928 9392 275980 9444
rect 281080 9392 281132 9444
rect 282828 9392 282880 9444
rect 283288 9392 283340 9444
rect 285404 9392 285456 9444
rect 289728 9392 289780 9444
rect 291016 9392 291068 9444
rect 292120 9392 292172 9444
rect 292948 9392 293000 9444
rect 294328 9392 294380 9444
rect 295524 9392 295576 9444
rect 300768 9392 300820 9444
rect 301872 9392 301924 9444
rect 302056 9392 302108 9444
rect 303160 9392 303212 9444
rect 309784 9392 309836 9444
rect 311532 9392 311584 9444
rect 324044 9392 324096 9444
rect 325056 9392 325108 9444
rect 326344 9392 326396 9444
rect 327080 9392 327132 9444
rect 328368 9392 328420 9444
rect 329656 9392 329708 9444
rect 340604 9392 340656 9444
rect 342168 9392 342220 9444
rect 349528 9392 349580 9444
rect 351828 9392 351880 9444
rect 352840 9392 352892 9444
rect 354496 9392 354548 9444
rect 358360 9392 358412 9444
rect 360108 9392 360160 9444
rect 361488 9392 361540 9444
rect 362868 9392 362920 9444
rect 367008 9392 367060 9444
rect 368296 9392 368348 9444
rect 369400 9392 369452 9444
rect 371148 9392 371200 9444
rect 374920 9392 374972 9444
rect 375380 9392 375432 9444
rect 390376 9392 390428 9444
rect 391848 9392 391900 9444
rect 401324 9392 401376 9444
rect 402888 9392 402940 9444
rect 405648 9392 405700 9444
rect 407028 9392 407080 9444
rect 410984 9392 411036 9444
rect 412548 9392 412600 9444
rect 414664 9392 414716 9444
rect 416688 9392 416740 9444
rect 417976 9392 418028 9444
rect 419448 9392 419500 9444
rect 432328 9392 432380 9444
rect 433340 9392 433392 9444
rect 437848 9392 437900 9444
rect 438860 9392 438912 9444
rect 443368 9392 443420 9444
rect 456892 9392 456944 9444
rect 457720 9392 457772 9444
rect 471888 9392 471940 9444
rect 473176 9392 473228 9444
rect 486332 9392 486384 9444
rect 489644 9392 489696 9444
rect 503628 9392 503680 9444
rect 505008 9392 505060 9444
rect 517612 9392 517664 9444
rect 522856 9392 522908 9444
rect 536012 9392 536064 9444
rect 34888 9324 34940 9376
rect 43076 9324 43128 9376
rect 43352 9324 43404 9376
rect 49700 9324 49752 9376
rect 50988 9324 51040 9376
rect 56600 9324 56652 9376
rect 64972 9324 65024 9376
rect 70676 9324 70728 9376
rect 81532 9324 81584 9376
rect 86132 9324 86184 9376
rect 95332 9324 95384 9376
rect 99380 9324 99432 9376
rect 133880 9324 133932 9376
rect 135812 9324 135864 9376
rect 143540 9324 143592 9376
rect 144920 9324 144972 9376
rect 282184 9324 282236 9376
rect 284208 9324 284260 9376
rect 316408 9324 316460 9376
rect 317420 9324 317472 9376
rect 320824 9324 320876 9376
rect 322848 9324 322900 9376
rect 331864 9324 331916 9376
rect 333888 9324 333940 9376
rect 337384 9324 337436 9376
rect 339408 9324 339460 9376
rect 377864 9324 377916 9376
rect 379428 9324 379480 9376
rect 387064 9324 387116 9376
rect 389088 9324 389140 9376
rect 393688 9324 393740 9376
rect 394792 9324 394844 9376
rect 398104 9324 398156 9376
rect 400128 9324 400180 9376
rect 433248 9324 433300 9376
rect 446220 9324 446272 9376
rect 456524 9324 456576 9376
rect 470508 9324 470560 9376
rect 476488 9324 476540 9376
rect 490104 9324 490156 9376
rect 496360 9324 496412 9376
rect 510160 9324 510212 9376
rect 514024 9324 514076 9376
rect 527916 9324 527968 9376
rect 529480 9324 529532 9376
rect 542360 9324 542412 9376
rect 23296 9256 23348 9308
rect 29000 9256 29052 9308
rect 29920 9256 29972 9308
rect 37556 9256 37608 9308
rect 46940 9256 46992 9308
rect 54116 9256 54168 9308
rect 56692 9256 56744 9308
rect 62948 9256 63000 9308
rect 63500 9256 63552 9308
rect 69572 9256 69624 9308
rect 70952 9256 71004 9308
rect 76196 9256 76248 9308
rect 79968 9256 80020 9308
rect 84200 9256 84252 9308
rect 304264 9256 304316 9308
rect 305736 9256 305788 9308
rect 342904 9256 342956 9308
rect 343732 9256 343784 9308
rect 359464 9256 359516 9308
rect 361488 9256 361540 9308
rect 403624 9256 403676 9308
rect 404360 9256 404412 9308
rect 415768 9256 415820 9308
rect 417976 9256 418028 9308
rect 429016 9256 429068 9308
rect 429660 9256 429712 9308
rect 436744 9256 436796 9308
rect 438676 9256 438728 9308
rect 438768 9256 438820 9308
rect 452108 9256 452160 9308
rect 455328 9256 455380 9308
rect 467840 9256 467892 9308
rect 482008 9256 482060 9308
rect 495532 9256 495584 9308
rect 504088 9256 504140 9308
rect 517520 9256 517572 9308
rect 519544 9256 519596 9308
rect 533988 9256 534040 9308
rect 538128 9256 538180 9308
rect 551836 9256 551888 9308
rect 25044 9188 25096 9240
rect 33140 9188 33192 9240
rect 44364 9188 44416 9240
rect 51908 9188 51960 9240
rect 53932 9188 53984 9240
rect 60740 9188 60792 9240
rect 72424 9188 72476 9240
rect 77300 9188 77352 9240
rect 92572 9188 92624 9240
rect 96068 9188 96120 9240
rect 199108 9188 199160 9240
rect 202052 9188 202104 9240
rect 275560 9188 275612 9240
rect 277124 9188 277176 9240
rect 332968 9188 333020 9240
rect 335084 9188 335136 9240
rect 344928 9188 344980 9240
rect 345112 9188 345164 9240
rect 382648 9188 382700 9240
rect 384396 9188 384448 9240
rect 442264 9188 442316 9240
rect 455696 9188 455748 9240
rect 458824 9188 458876 9240
rect 471980 9188 472032 9240
rect 475384 9188 475436 9240
rect 488540 9188 488592 9240
rect 490840 9188 490892 9240
rect 505008 9188 505060 9240
rect 507400 9188 507452 9240
rect 520464 9188 520516 9240
rect 525064 9188 525116 9240
rect 538864 9188 538916 9240
rect 17868 9120 17920 9172
rect 18788 9120 18840 9172
rect 24032 9120 24084 9172
rect 32036 9120 32088 9172
rect 32772 9120 32824 9172
rect 40040 9120 40092 9172
rect 41512 9120 41564 9172
rect 48596 9120 48648 9172
rect 49608 9120 49660 9172
rect 55312 9120 55364 9172
rect 62672 9120 62724 9172
rect 68468 9120 68520 9172
rect 87788 9120 87840 9172
rect 91652 9120 91704 9172
rect 92480 9120 92532 9172
rect 97172 9120 97224 9172
rect 111984 9120 112036 9172
rect 114836 9120 114888 9172
rect 201500 9120 201552 9172
rect 204260 9120 204312 9172
rect 210976 9120 211028 9172
rect 213092 9120 213144 9172
rect 263416 9120 263468 9172
rect 264152 9120 264204 9172
rect 268936 9120 268988 9172
rect 270040 9120 270092 9172
rect 298744 9120 298796 9172
rect 300676 9120 300728 9172
rect 318616 9120 318668 9172
rect 320088 9120 320140 9172
rect 329564 9120 329616 9172
rect 331128 9120 331180 9172
rect 425704 9120 425756 9172
rect 427728 9120 427780 9172
rect 440056 9120 440108 9172
rect 453304 9120 453356 9172
rect 23388 9052 23440 9104
rect 30932 9052 30984 9104
rect 31668 9052 31720 9104
rect 38660 9052 38712 9104
rect 82820 9052 82872 9104
rect 87236 9052 87288 9104
rect 90180 9052 90232 9104
rect 93952 9052 94004 9104
rect 373724 9052 373776 9104
rect 374368 9052 374420 9104
rect 377128 9052 377180 9104
rect 379244 9052 379296 9104
rect 427544 9052 427596 9104
rect 440332 9052 440384 9104
rect 447784 9052 447836 9104
rect 37280 8984 37332 9036
rect 45560 8984 45612 9036
rect 73160 8984 73212 9036
rect 78680 8984 78732 9036
rect 97172 8984 97224 9036
rect 100760 8984 100812 9036
rect 102140 8984 102192 9036
rect 106280 8984 106332 9036
rect 118056 8984 118108 9036
rect 120356 8984 120408 9036
rect 212172 8984 212224 9036
rect 214196 8984 214248 9036
rect 362776 8984 362828 9036
rect 363328 8984 363380 9036
rect 364984 8984 365036 9036
rect 365720 8984 365772 9036
rect 371608 8984 371660 9036
rect 372620 8984 372672 9036
rect 435640 8984 435692 9036
rect 448612 8984 448664 9036
rect 449808 9052 449860 9104
rect 462320 9120 462372 9172
rect 465448 9120 465500 9172
rect 480168 9120 480220 9172
rect 480904 9120 480956 9172
rect 495348 9120 495400 9172
rect 497464 9120 497516 9172
rect 510712 9120 510764 9172
rect 517336 9120 517388 9172
rect 530032 9120 530084 9172
rect 541624 9120 541676 9172
rect 555424 9120 555476 9172
rect 464344 9052 464396 9104
rect 478788 9052 478840 9104
rect 484216 9052 484268 9104
rect 496912 9052 496964 9104
rect 500776 9052 500828 9104
rect 514668 9052 514720 9104
rect 523960 9052 524012 9104
rect 538036 9052 538088 9104
rect 544936 9052 544988 9104
rect 557632 9052 557684 9104
rect 461584 8984 461636 9036
rect 462136 8984 462188 9036
rect 475108 8984 475160 9036
rect 477408 8984 477460 9036
rect 490012 8984 490064 9036
rect 493048 8984 493100 9036
rect 506480 8984 506532 9036
rect 520648 8984 520700 9036
rect 534908 8984 534960 9036
rect 537208 8984 537260 9036
rect 551928 8984 551980 9036
rect 15200 8916 15252 8968
rect 20996 8916 21048 8968
rect 27620 8916 27672 8968
rect 36452 8916 36504 8968
rect 43444 8916 43496 8968
rect 51080 8916 51132 8968
rect 53104 8916 53156 8968
rect 59636 8916 59688 8968
rect 60924 8916 60976 8968
rect 67640 8916 67692 8968
rect 353944 8916 353996 8968
rect 355048 8916 355100 8968
rect 402520 8916 402572 8968
rect 403440 8916 403492 8968
rect 431224 8916 431276 8968
rect 432236 8916 432288 8968
rect 434536 8916 434588 8968
rect 447416 8916 447468 8968
rect 451096 8916 451148 8968
rect 464988 8916 465040 8968
rect 470968 8916 471020 8968
rect 484676 8916 484728 8968
rect 487528 8916 487580 8968
rect 500960 8916 501012 8968
rect 510528 8916 510580 8968
rect 524236 8916 524288 8968
rect 530584 8916 530636 8968
rect 545028 8916 545080 8968
rect 547972 8916 548024 8968
rect 568488 8916 568540 8968
rect 22100 8848 22152 8900
rect 25412 8848 25464 8900
rect 55220 8848 55272 8900
rect 62120 8848 62172 8900
rect 85580 8848 85632 8900
rect 90548 8848 90600 8900
rect 126520 8848 126572 8900
rect 128360 8848 128412 8900
rect 265624 8848 265676 8900
rect 266544 8848 266596 8900
rect 285496 8848 285548 8900
rect 286048 8848 286100 8900
rect 288808 8848 288860 8900
rect 291108 8848 291160 8900
rect 313096 8848 313148 8900
rect 314568 8848 314620 8900
rect 360568 8848 360620 8900
rect 362776 8848 362828 8900
rect 388168 8848 388220 8900
rect 390192 8848 390244 8900
rect 399208 8848 399260 8900
rect 401508 8848 401560 8900
rect 471704 8848 471756 8900
rect 485688 8848 485740 8900
rect 488448 8848 488500 8900
rect 501052 8848 501104 8900
rect 506296 8848 506348 8900
rect 518900 8848 518952 8900
rect 521568 8848 521620 8900
rect 535368 8848 535420 8900
rect 363880 8780 363932 8832
rect 364800 8780 364852 8832
rect 446680 8780 446732 8832
rect 460388 8780 460440 8832
rect 460848 8780 460900 8832
rect 474648 8780 474700 8832
rect 479800 8780 479852 8832
rect 493968 8780 494020 8832
rect 508504 8780 508556 8832
rect 522948 8780 523000 8832
rect 531504 8780 531556 8832
rect 545764 8780 545816 8832
rect 108212 8712 108264 8764
rect 110420 8712 110472 8764
rect 223948 8712 224000 8764
rect 225236 8712 225288 8764
rect 231032 8712 231084 8764
rect 231860 8712 231912 8764
rect 404728 8712 404780 8764
rect 406108 8712 406160 8764
rect 420184 8712 420236 8764
rect 420920 8712 420972 8764
rect 453212 8712 453264 8764
rect 467472 8712 467524 8764
rect 474280 8712 474332 8764
rect 487160 8712 487212 8764
rect 495256 8712 495308 8764
rect 507860 8712 507912 8764
rect 511816 8712 511868 8764
rect 525708 8712 525760 8764
rect 525800 8712 525852 8764
rect 539692 8712 539744 8764
rect 344008 8644 344060 8696
rect 345020 8644 345072 8696
rect 452200 8644 452252 8696
rect 466276 8644 466328 8696
rect 468760 8644 468812 8696
rect 481640 8644 481692 8696
rect 485320 8644 485372 8696
rect 498200 8644 498252 8696
rect 512920 8644 512972 8696
rect 526444 8644 526496 8696
rect 84292 8576 84344 8628
rect 89720 8576 89772 8628
rect 348424 8576 348476 8628
rect 350448 8576 350500 8628
rect 368204 8576 368256 8628
rect 369768 8576 369820 8628
rect 424600 8576 424652 8628
rect 426072 8576 426124 8628
rect 441160 8576 441212 8628
rect 454500 8576 454552 8628
rect 466368 8576 466420 8628
rect 478880 8576 478932 8628
rect 491944 8576 491996 8628
rect 505560 8576 505612 8628
rect 515128 8576 515180 8628
rect 528560 8576 528612 8628
rect 267648 8508 267700 8560
rect 268844 8508 268896 8560
rect 306288 8508 306340 8560
rect 306472 8508 306524 8560
rect 315304 8508 315356 8560
rect 316040 8508 316092 8560
rect 383568 8508 383620 8560
rect 383660 8508 383712 8560
rect 392584 8508 392636 8560
rect 393320 8508 393372 8560
rect 421288 8508 421340 8560
rect 423036 8508 423088 8560
rect 430120 8508 430172 8560
rect 430948 8508 431000 8560
rect 454408 8508 454460 8560
rect 468668 8508 468720 8560
rect 498568 8508 498620 8560
rect 513288 8508 513340 8560
rect 207388 8440 207440 8492
rect 209872 8440 209924 8492
rect 229836 8440 229888 8492
rect 230756 8440 230808 8492
rect 310888 8440 310940 8492
rect 312728 8440 312780 8492
rect 459928 8440 459980 8492
rect 474556 8440 474608 8492
rect 493784 8440 493836 8492
rect 506756 8440 506808 8492
rect 509608 8440 509660 8492
rect 524328 8440 524380 8492
rect 60556 8372 60608 8424
rect 65156 8372 65208 8424
rect 69940 8372 69992 8424
rect 75092 8372 75144 8424
rect 100944 8372 100996 8424
rect 103796 8372 103848 8424
rect 208584 8372 208636 8424
rect 211160 8372 211212 8424
rect 219256 8372 219308 8424
rect 220820 8372 220872 8424
rect 232228 8372 232280 8424
rect 233240 8372 233292 8424
rect 257896 8372 257948 8424
rect 258264 8372 258316 8424
rect 276664 8372 276716 8424
rect 278320 8372 278372 8424
rect 379336 8372 379388 8424
rect 380808 8372 380860 8424
rect 412456 8372 412508 8424
rect 412640 8372 412692 8424
rect 13820 8304 13872 8356
rect 16672 8304 16724 8356
rect 16764 8304 16816 8356
rect 19892 8304 19944 8356
rect 39304 8304 39356 8356
rect 46388 8304 46440 8356
rect 52092 8304 52144 8356
rect 57428 8304 57480 8356
rect 60004 8304 60056 8356
rect 66260 8304 66312 8356
rect 80520 8304 80572 8356
rect 85028 8304 85080 8356
rect 91192 8304 91244 8356
rect 95240 8304 95292 8356
rect 100852 8304 100904 8356
rect 104900 8304 104952 8356
rect 110512 8304 110564 8356
rect 113732 8304 113784 8356
rect 120172 8304 120224 8356
rect 122932 8304 122984 8356
rect 197912 8304 197964 8356
rect 200948 8304 201000 8356
rect 218060 8304 218112 8356
rect 219716 8304 219768 8356
rect 238116 8304 238168 8356
rect 238760 8304 238812 8356
rect 266728 8304 266780 8356
rect 267740 8304 267792 8356
rect 286600 8304 286652 8356
rect 287244 8304 287296 8356
rect 296536 8304 296588 8356
rect 296720 8304 296772 8356
rect 305368 8304 305420 8356
rect 306932 8304 306984 8356
rect 335176 8304 335228 8356
rect 335360 8304 335412 8356
rect 422208 8304 422260 8356
rect 422300 8304 422352 8356
rect 3424 6468 3476 6520
rect 8944 6468 8996 6520
rect 5264 4088 5316 4140
rect 15200 4088 15252 4140
rect 30104 4088 30156 4140
rect 35992 4088 36044 4140
rect 39580 4088 39632 4140
rect 45744 4088 45796 4140
rect 50160 4088 50212 4140
rect 56692 4088 56744 4140
rect 58440 4088 58492 4140
rect 64972 4088 65024 4140
rect 67916 4088 67968 4140
rect 74632 4088 74684 4140
rect 79692 4088 79744 4140
rect 85580 4088 85632 4140
rect 89168 4088 89220 4140
rect 95240 4088 95292 4140
rect 97448 4088 97500 4140
rect 103612 4088 103664 4140
rect 108120 4088 108172 4140
rect 114560 4088 114612 4140
rect 116400 4088 116452 4140
rect 124128 4088 124180 4140
rect 128176 4088 128228 4140
rect 133880 4088 133932 4140
rect 137652 4088 137704 4140
rect 143540 4088 143592 4140
rect 145932 4088 145984 4140
rect 151820 4088 151872 4140
rect 157800 4088 157852 4140
rect 162860 4088 162912 4140
rect 296260 4088 296312 4140
rect 298468 4088 298520 4140
rect 324228 4088 324280 4140
rect 326804 4088 326856 4140
rect 333888 4088 333940 4140
rect 337476 4088 337528 4140
rect 342168 4088 342220 4140
rect 346952 4088 347004 4140
rect 351828 4088 351880 4140
rect 356336 4088 356388 4140
rect 358728 4088 358780 4140
rect 364616 4088 364668 4140
rect 368296 4088 368348 4140
rect 375288 4088 375340 4140
rect 387708 4088 387760 4140
rect 395344 4088 395396 4140
rect 416688 4088 416740 4140
rect 426164 4088 426216 4140
rect 506756 4088 506808 4140
rect 511264 4088 511316 4140
rect 516508 4088 516560 4140
rect 520740 4088 520792 4140
rect 525708 4088 525760 4140
rect 530124 4088 530176 4140
rect 535368 4088 535420 4140
rect 540796 4088 540848 4140
rect 542728 4088 542780 4140
rect 563244 4088 563296 4140
rect 14740 4020 14792 4072
rect 24952 4020 25004 4072
rect 53748 4020 53800 4072
rect 60004 4020 60056 4072
rect 62028 4020 62080 4072
rect 68652 4020 68704 4072
rect 69112 4020 69164 4072
rect 76104 4020 76156 4072
rect 77392 4020 77444 4072
rect 84384 4020 84436 4072
rect 125876 4020 125928 4072
rect 133788 4020 133840 4072
rect 136456 4020 136508 4072
rect 143448 4020 143500 4072
rect 155408 4020 155460 4072
rect 161572 4020 161624 4072
rect 177856 4020 177908 4072
rect 182180 4020 182232 4072
rect 187332 4020 187384 4072
rect 190460 4020 190512 4072
rect 196808 4020 196860 4072
rect 200212 4020 200264 4072
rect 340696 4020 340748 4072
rect 345756 4020 345808 4072
rect 350448 4020 350500 4072
rect 355232 4020 355284 4072
rect 361488 4020 361540 4072
rect 367008 4020 367060 4072
rect 369768 4020 369820 4072
rect 376484 4020 376536 4072
rect 406108 4020 406160 4072
rect 415492 4020 415544 4072
rect 423036 4020 423088 4072
rect 433248 4020 433300 4072
rect 524236 4020 524288 4072
rect 529020 4020 529072 4072
rect 539416 4020 539468 4072
rect 559748 4020 559800 4072
rect 9956 3952 10008 4004
rect 22100 3952 22152 4004
rect 24216 3952 24268 4004
rect 31668 3952 31720 4004
rect 54944 3952 54996 4004
rect 60924 3952 60976 4004
rect 111616 3952 111668 4004
rect 118056 3952 118108 4004
rect 118792 3952 118844 4004
rect 126888 3952 126940 4004
rect 166080 3952 166132 4004
rect 171140 3952 171192 4004
rect 313188 3952 313240 4004
rect 316224 3952 316276 4004
rect 324136 3952 324188 4004
rect 328000 3952 328052 4004
rect 360108 3952 360160 4004
rect 365812 3952 365864 4004
rect 378048 3952 378100 4004
rect 384764 3952 384816 4004
rect 389088 3952 389140 4004
rect 396540 3952 396592 4004
rect 401508 3952 401560 4004
rect 409604 3952 409656 4004
rect 412364 3952 412416 4004
rect 421380 3952 421432 4004
rect 422300 3952 422352 4004
rect 434444 3952 434496 4004
rect 488540 3952 488592 4004
rect 491116 3952 491168 4004
rect 498200 3952 498252 4004
rect 501788 3952 501840 4004
rect 533988 3952 534040 4004
rect 538404 3952 538456 4004
rect 540520 3952 540572 4004
rect 560852 3952 560904 4004
rect 4068 3884 4120 3936
rect 16672 3884 16724 3936
rect 18052 3884 18104 3936
rect 23664 3884 23716 3936
rect 44272 3884 44324 3936
rect 52092 3884 52144 3936
rect 101036 3884 101088 3936
rect 108212 3884 108264 3936
rect 332508 3884 332560 3936
rect 336280 3884 336332 3936
rect 372620 3884 372672 3936
rect 379980 3884 380032 3936
rect 392492 3884 392544 3936
rect 401324 3884 401376 3936
rect 401416 3884 401468 3936
rect 410800 3884 410852 3936
rect 411168 3884 411220 3936
rect 420184 3884 420236 3936
rect 427728 3884 427780 3936
rect 437940 3884 437992 3936
rect 534908 3884 534960 3936
rect 539600 3884 539652 3936
rect 545028 3884 545080 3936
rect 550272 3884 550324 3936
rect 552020 3884 552072 3936
rect 553216 3884 553268 3936
rect 553400 3884 553452 3936
rect 575112 3884 575164 3936
rect 2872 3816 2924 3868
rect 17868 3816 17920 3868
rect 21824 3816 21876 3868
rect 27620 3816 27672 3868
rect 31300 3816 31352 3868
rect 37280 3816 37332 3868
rect 71504 3816 71556 3868
rect 78588 3816 78640 3868
rect 80888 3816 80940 3868
rect 87788 3816 87840 3868
rect 122288 3816 122340 3868
rect 129648 3816 129700 3868
rect 141240 3816 141292 3868
rect 147680 3816 147732 3868
rect 150624 3816 150676 3868
rect 155960 3816 156012 3868
rect 167184 3816 167236 3868
rect 172612 3816 172664 3868
rect 188528 3816 188580 3868
rect 191932 3816 191984 3868
rect 286048 3816 286100 3868
rect 287796 3816 287848 3868
rect 295524 3816 295576 3868
rect 297272 3816 297324 3868
rect 305736 3816 305788 3868
rect 307944 3816 307996 3868
rect 315856 3816 315908 3868
rect 318524 3816 318576 3868
rect 362776 3816 362828 3868
rect 368204 3816 368256 3868
rect 394792 3816 394844 3868
rect 403624 3816 403676 3868
rect 407396 3816 407448 3868
rect 417884 3816 417936 3868
rect 418068 3816 418120 3868
rect 428464 3816 428516 3868
rect 429660 3816 429712 3868
rect 441528 3816 441580 3868
rect 536012 3816 536064 3868
rect 541992 3816 542044 3868
rect 542360 3816 542412 3868
rect 549076 3816 549128 3868
rect 553492 3816 553544 3868
rect 576308 3816 576360 3868
rect 572 3748 624 3800
rect 13820 3748 13872 3800
rect 15936 3748 15988 3800
rect 23388 3748 23440 3800
rect 25320 3748 25372 3800
rect 32772 3748 32824 3800
rect 34796 3748 34848 3800
rect 41512 3748 41564 3800
rect 43076 3748 43128 3800
rect 50988 3748 51040 3800
rect 51356 3748 51408 3800
rect 59268 3748 59320 3800
rect 64328 3748 64380 3800
rect 70952 3748 71004 3800
rect 99840 3748 99892 3800
rect 106832 3748 106884 3800
rect 163688 3748 163740 3800
rect 168380 3748 168432 3800
rect 335176 3748 335228 3800
rect 338672 3748 338724 3800
rect 362868 3748 362920 3800
rect 369400 3748 369452 3800
rect 372160 3748 372212 3800
rect 378876 3748 378928 3800
rect 379428 3748 379480 3800
rect 387156 3748 387208 3800
rect 391848 3748 391900 3800
rect 400036 3748 400088 3800
rect 400128 3748 400180 3800
rect 408408 3748 408460 3800
rect 420828 3748 420880 3800
rect 430856 3748 430908 3800
rect 430948 3748 431000 3800
rect 442632 3748 442684 3800
rect 478880 3748 478932 3800
rect 481732 3748 481784 3800
rect 538036 3748 538088 3800
rect 543188 3748 543240 3800
rect 550640 3748 550692 3800
rect 552756 3748 552808 3800
rect 554780 3748 554832 3800
rect 577412 3748 577464 3800
rect 11152 3680 11204 3732
rect 26240 3680 26292 3732
rect 32404 3680 32456 3732
rect 39304 3680 39356 3732
rect 41880 3680 41932 3732
rect 49608 3680 49660 3732
rect 73804 3680 73856 3732
rect 80520 3680 80572 3732
rect 92756 3680 92808 3732
rect 99472 3680 99524 3732
rect 106924 3680 106976 3732
rect 113272 3680 113324 3732
rect 121092 3680 121144 3732
rect 128268 3680 128320 3732
rect 140044 3680 140096 3732
rect 146300 3680 146352 3732
rect 148324 3680 148376 3732
rect 154580 3680 154632 3732
rect 160100 3680 160152 3732
rect 165620 3680 165672 3732
rect 171968 3680 172020 3732
rect 176660 3680 176712 3732
rect 304448 3680 304500 3732
rect 306748 3680 306800 3732
rect 354496 3680 354548 3732
rect 359924 3680 359976 3732
rect 382924 3680 382976 3732
rect 390652 3680 390704 3732
rect 394884 3680 394936 3732
rect 404820 3680 404872 3732
rect 407028 3680 407080 3732
rect 416688 3680 416740 3732
rect 423772 3680 423824 3732
rect 435548 3680 435600 3732
rect 438676 3680 438728 3732
rect 449808 3680 449860 3732
rect 527916 3680 527968 3732
rect 532516 3680 532568 3732
rect 545764 3680 545816 3732
rect 551468 3680 551520 3732
rect 556160 3680 556212 3732
rect 578608 3680 578660 3732
rect 6460 3612 6512 3664
rect 22192 3612 22244 3664
rect 23020 3612 23072 3664
rect 29920 3612 29972 3664
rect 63224 3612 63276 3664
rect 69940 3612 69992 3664
rect 72608 3612 72660 3664
rect 79968 3612 80020 3664
rect 104532 3612 104584 3664
rect 110512 3612 110564 3664
rect 130568 3612 130620 3664
rect 137928 3612 137980 3664
rect 138848 3612 138900 3664
rect 145104 3612 145156 3664
rect 158904 3612 158956 3664
rect 164240 3612 164292 3664
rect 169576 3612 169628 3664
rect 173900 3612 173952 3664
rect 353208 3612 353260 3664
rect 358728 3612 358780 3664
rect 363328 3612 363380 3664
rect 370596 3612 370648 3664
rect 371148 3612 371200 3664
rect 377680 3612 377732 3664
rect 385040 3612 385092 3664
rect 12348 3544 12400 3596
rect 27804 3544 27856 3596
rect 33600 3544 33652 3596
rect 41328 3544 41380 3596
rect 59636 3544 59688 3596
rect 66352 3544 66404 3596
rect 82084 3544 82136 3596
rect 89628 3544 89680 3596
rect 90364 3544 90416 3596
rect 97172 3544 97224 3596
rect 109316 3544 109368 3596
rect 117228 3544 117280 3596
rect 131764 3544 131816 3596
rect 139308 3544 139360 3596
rect 170772 3544 170824 3596
rect 175280 3544 175332 3596
rect 180248 3544 180300 3596
rect 183652 3544 183704 3596
rect 259460 3544 259512 3596
rect 260656 3544 260708 3596
rect 303160 3544 303212 3596
rect 305552 3544 305604 3596
rect 346400 3544 346452 3596
rect 352840 3544 352892 3596
rect 368388 3544 368440 3596
rect 374092 3544 374144 3596
rect 380808 3544 380860 3596
rect 388260 3544 388312 3596
rect 402888 3612 402940 3664
rect 411904 3612 411956 3664
rect 412548 3612 412600 3664
rect 422576 3612 422628 3664
rect 427820 3612 427872 3664
rect 439136 3612 439188 3664
rect 551836 3612 551888 3664
rect 558552 3612 558604 3664
rect 560300 3612 560352 3664
rect 583392 3612 583444 3664
rect 394240 3544 394292 3596
rect 396264 3544 396316 3596
rect 7656 3476 7708 3528
rect 18052 3476 18104 3528
rect 18236 3476 18288 3528
rect 25044 3476 25096 3528
rect 26516 3476 26568 3528
rect 33784 3476 33836 3528
rect 37188 3476 37240 3528
rect 43444 3476 43496 3528
rect 47860 3476 47912 3528
rect 53932 3476 53984 3528
rect 57244 3476 57296 3528
rect 63500 3476 63552 3528
rect 75000 3476 75052 3528
rect 81532 3476 81584 3528
rect 83280 3476 83332 3528
rect 90180 3476 90232 3528
rect 91560 3476 91612 3528
rect 98460 3476 98512 3528
rect 103336 3476 103388 3528
rect 109132 3476 109184 3528
rect 112812 3476 112864 3528
rect 118700 3476 118752 3528
rect 151820 3476 151872 3528
rect 157340 3476 157392 3528
rect 168380 3476 168432 3528
rect 172520 3476 172572 3528
rect 174268 3476 174320 3528
rect 178132 3476 178184 3528
rect 179052 3476 179104 3528
rect 183560 3476 183612 3528
rect 183744 3476 183796 3528
rect 187700 3476 187752 3528
rect 189724 3476 189776 3528
rect 193312 3476 193364 3528
rect 291016 3476 291068 3528
rect 292580 3476 292632 3528
rect 292948 3476 293000 3528
rect 294880 3476 294932 3528
rect 300676 3476 300728 3528
rect 301964 3476 302016 3528
rect 306932 3476 306984 3528
rect 309048 3476 309100 3528
rect 310428 3476 310480 3528
rect 312636 3476 312688 3528
rect 316040 3476 316092 3528
rect 319720 3476 319772 3528
rect 322848 3476 322900 3528
rect 325608 3476 325660 3528
rect 329748 3476 329800 3528
rect 332692 3476 332744 3528
rect 334256 3476 334308 3528
rect 339868 3476 339920 3528
rect 343548 3476 343600 3528
rect 348056 3476 348108 3528
rect 355048 3476 355100 3528
rect 361120 3476 361172 3528
rect 390468 3476 390520 3528
rect 398932 3476 398984 3528
rect 403440 3544 403492 3596
rect 413100 3544 413152 3596
rect 420920 3544 420972 3596
rect 432052 3544 432104 3596
rect 432236 3544 432288 3596
rect 443828 3544 443880 3596
rect 471980 3544 472032 3596
rect 473452 3544 473504 3596
rect 491392 3544 491444 3596
rect 494704 3544 494756 3596
rect 507860 3544 507912 3596
rect 512460 3544 512512 3596
rect 516048 3544 516100 3596
rect 519544 3544 519596 3596
rect 526444 3544 526496 3596
rect 531320 3544 531372 3596
rect 531412 3544 531464 3596
rect 406016 3476 406068 3528
rect 412640 3476 412692 3528
rect 423772 3476 423824 3528
rect 426072 3476 426124 3528
rect 436744 3476 436796 3528
rect 438860 3476 438912 3528
rect 450912 3476 450964 3528
rect 462320 3476 462372 3528
rect 463976 3476 464028 3528
rect 467840 3476 467892 3528
rect 469864 3476 469916 3528
rect 474648 3476 474700 3528
rect 475752 3476 475804 3528
rect 476304 3476 476356 3528
rect 478144 3476 478196 3528
rect 480628 3476 480680 3528
rect 482836 3476 482888 3528
rect 484308 3476 484360 3528
rect 485228 3476 485280 3528
rect 490104 3476 490156 3528
rect 492312 3476 492364 3528
rect 496452 3476 496504 3528
rect 499396 3476 499448 3528
rect 499672 3476 499724 3528
rect 502984 3476 503036 3528
rect 505560 3476 505612 3528
rect 508872 3476 508924 3528
rect 513288 3476 513340 3528
rect 515956 3476 516008 3528
rect 517520 3476 517572 3528
rect 521844 3476 521896 3528
rect 524328 3476 524380 3528
rect 527824 3476 527876 3528
rect 528560 3476 528612 3528
rect 533712 3476 533764 3528
rect 538864 3544 538916 3596
rect 544384 3544 544436 3596
rect 547880 3544 547932 3596
rect 554964 3544 555016 3596
rect 558920 3544 558972 3596
rect 581000 3544 581052 3596
rect 1676 3408 1728 3460
rect 18144 3408 18196 3460
rect 19432 3408 19484 3460
rect 26424 3408 26476 3460
rect 45468 3408 45520 3460
rect 52276 3408 52328 3460
rect 52552 3408 52604 3460
rect 60556 3408 60608 3460
rect 60832 3408 60884 3460
rect 68928 3408 68980 3460
rect 70308 3408 70360 3460
rect 75920 3408 75972 3460
rect 85672 3408 85724 3460
rect 92572 3408 92624 3460
rect 95148 3408 95200 3460
rect 100852 3408 100904 3460
rect 102232 3408 102284 3460
rect 109224 3408 109276 3460
rect 110512 3408 110564 3460
rect 118608 3408 118660 3460
rect 119896 3408 119948 3460
rect 126520 3408 126572 3460
rect 129372 3408 129424 3460
rect 136548 3408 136600 3460
rect 142436 3408 142488 3460
rect 149060 3408 149112 3460
rect 149520 3408 149572 3460
rect 156052 3408 156104 3460
rect 161296 3408 161348 3460
rect 167092 3408 167144 3460
rect 175464 3408 175516 3460
rect 179420 3408 179472 3460
rect 181444 3408 181496 3460
rect 184940 3408 184992 3460
rect 190828 3408 190880 3460
rect 194784 3408 194836 3460
rect 301320 3408 301372 3460
rect 303160 3408 303212 3460
rect 307760 3408 307812 3460
rect 311440 3408 311492 3460
rect 311532 3408 311584 3460
rect 313832 3408 313884 3460
rect 317512 3408 317564 3460
rect 322112 3408 322164 3460
rect 325056 3408 325108 3460
rect 329196 3408 329248 3460
rect 329656 3408 329708 3460
rect 333888 3408 333940 3460
rect 343732 3408 343784 3460
rect 349252 3408 349304 3460
rect 351092 3408 351144 3460
rect 357532 3408 357584 3460
rect 365720 3408 365772 3460
rect 372896 3408 372948 3460
rect 373356 3408 373408 3460
rect 381176 3408 381228 3460
rect 381728 3408 381780 3460
rect 389456 3408 389508 3460
rect 390192 3408 390244 3460
rect 397736 3408 397788 3460
rect 398748 3408 398800 3460
rect 407212 3408 407264 3460
rect 414020 3408 414072 3460
rect 13544 3340 13596 3392
rect 23296 3340 23348 3392
rect 27712 3340 27764 3392
rect 34704 3340 34756 3392
rect 65524 3340 65576 3392
rect 72424 3340 72476 3392
rect 96252 3340 96304 3392
rect 102140 3340 102192 3392
rect 115204 3340 115256 3392
rect 122748 3340 122800 3392
rect 301872 3340 301924 3392
rect 304356 3340 304408 3392
rect 335360 3340 335412 3392
rect 340972 3340 341024 3392
rect 345112 3340 345164 3392
rect 351644 3340 351696 3392
rect 393320 3340 393372 3392
rect 402520 3340 402572 3392
rect 404360 3340 404412 3392
rect 414296 3340 414348 3392
rect 417976 3340 418028 3392
rect 419448 3408 419500 3460
rect 429660 3408 429712 3460
rect 433340 3408 433392 3460
rect 445024 3408 445076 3460
rect 481640 3408 481692 3460
rect 484032 3408 484084 3460
rect 487160 3408 487212 3460
rect 489920 3408 489972 3460
rect 501052 3408 501104 3460
rect 505376 3408 505428 3460
rect 506480 3408 506532 3460
rect 510068 3408 510120 3460
rect 510712 3408 510764 3460
rect 514760 3408 514812 3460
rect 517612 3408 517664 3460
rect 523040 3408 523092 3460
rect 532608 3408 532660 3460
rect 537208 3408 537260 3460
rect 551928 3476 551980 3528
rect 557356 3476 557408 3528
rect 552664 3408 552716 3460
rect 552756 3408 552808 3460
rect 572720 3476 572772 3528
rect 557540 3408 557592 3460
rect 579804 3408 579856 3460
rect 8760 3272 8812 3324
rect 17960 3272 18012 3324
rect 20628 3272 20680 3324
rect 26332 3272 26384 3324
rect 40684 3272 40736 3324
rect 46940 3272 46992 3324
rect 48964 3272 49016 3324
rect 55220 3272 55272 3324
rect 78588 3272 78640 3324
rect 84292 3272 84344 3324
rect 87972 3272 88024 3324
rect 93860 3272 93912 3324
rect 117596 3272 117648 3324
rect 124220 3272 124272 3324
rect 143540 3272 143592 3324
rect 150440 3272 150492 3324
rect 154212 3272 154264 3324
rect 160192 3272 160244 3324
rect 162492 3272 162544 3324
rect 167000 3272 167052 3324
rect 176660 3272 176712 3324
rect 180800 3272 180852 3324
rect 186136 3272 186188 3324
rect 189172 3272 189224 3324
rect 194416 3272 194468 3324
rect 197452 3272 197504 3324
rect 202696 3272 202748 3324
rect 205732 3272 205784 3324
rect 296720 3272 296772 3324
rect 299664 3272 299716 3324
rect 306472 3272 306524 3324
rect 310244 3272 310296 3324
rect 314568 3272 314620 3324
rect 317328 3272 317380 3324
rect 317420 3272 317472 3324
rect 320916 3272 320968 3324
rect 326252 3272 326304 3324
rect 330392 3272 330444 3324
rect 331128 3272 331180 3324
rect 335084 3272 335136 3324
rect 339408 3272 339460 3324
rect 343364 3272 343416 3324
rect 345020 3272 345072 3324
rect 350448 3272 350500 3324
rect 379336 3272 379388 3324
rect 385960 3272 386012 3324
rect 408500 3272 408552 3324
rect 418988 3272 419040 3324
rect 424968 3340 425020 3392
rect 513196 3340 513248 3392
rect 517152 3340 517204 3392
rect 520464 3340 520516 3392
rect 525432 3340 525484 3392
rect 530032 3340 530084 3392
rect 536104 3340 536156 3392
rect 545120 3340 545172 3392
rect 427268 3272 427320 3324
rect 500960 3272 501012 3324
rect 504180 3272 504232 3324
rect 510160 3272 510212 3324
rect 513564 3272 513616 3324
rect 135260 3204 135312 3256
rect 142160 3204 142212 3256
rect 164884 3204 164936 3256
rect 169760 3204 169812 3256
rect 184940 3204 184992 3256
rect 189080 3204 189132 3256
rect 195612 3204 195664 3256
rect 198832 3204 198884 3256
rect 320088 3204 320140 3256
rect 323308 3204 323360 3256
rect 340788 3204 340840 3256
rect 344560 3204 344612 3256
rect 356060 3204 356112 3256
rect 363512 3204 363564 3256
rect 503628 3204 503680 3256
rect 506480 3204 506532 3256
rect 518900 3204 518952 3256
rect 524236 3204 524288 3256
rect 540980 3204 541032 3256
rect 547880 3204 547932 3256
rect 557632 3340 557684 3392
rect 565636 3340 565688 3392
rect 553216 3272 553268 3324
rect 573916 3272 573968 3324
rect 566832 3204 566884 3256
rect 17040 3136 17092 3188
rect 24032 3136 24084 3188
rect 98644 3136 98696 3188
rect 104992 3136 105044 3188
rect 126980 3136 127032 3188
rect 133972 3136 134024 3188
rect 173164 3136 173216 3188
rect 178040 3136 178092 3188
rect 182548 3136 182600 3188
rect 186320 3136 186372 3188
rect 291660 3136 291712 3188
rect 293684 3136 293736 3188
rect 298100 3136 298152 3188
rect 300768 3136 300820 3188
rect 312728 3136 312780 3188
rect 315028 3136 315080 3188
rect 321468 3136 321520 3188
rect 324412 3136 324464 3188
rect 327080 3136 327132 3188
rect 331588 3136 331640 3188
rect 486332 3136 486384 3188
rect 488816 3136 488868 3188
rect 490012 3136 490064 3188
rect 493508 3136 493560 3188
rect 495532 3136 495584 3188
rect 498200 3136 498252 3188
rect 505008 3136 505060 3188
rect 507676 3136 507728 3188
rect 514668 3136 514720 3188
rect 518348 3136 518400 3188
rect 522948 3136 523000 3188
rect 526628 3136 526680 3188
rect 555424 3136 555476 3188
rect 562048 3136 562100 3188
rect 374368 3068 374420 3120
rect 382372 3068 382424 3120
rect 38384 3000 38436 3052
rect 44364 3000 44416 3052
rect 76196 3000 76248 3052
rect 82820 3000 82872 3052
rect 84476 3000 84528 3052
rect 91192 3000 91244 3052
rect 114008 3000 114060 3052
rect 120172 3000 120224 3052
rect 123484 3000 123536 3052
rect 131028 3000 131080 3052
rect 134156 3000 134208 3052
rect 140780 3000 140832 3052
rect 144736 3000 144788 3052
rect 150532 3000 150584 3052
rect 278780 3000 278832 3052
rect 280712 3000 280764 3052
rect 284668 3000 284720 3052
rect 286600 3000 286652 3052
rect 288440 3000 288492 3052
rect 290188 3000 290240 3052
rect 294236 3000 294288 3052
rect 296076 3000 296128 3052
rect 356152 3000 356204 3052
rect 362316 3000 362368 3052
rect 364800 3000 364852 3052
rect 371700 3000 371752 3052
rect 383660 3000 383712 3052
rect 393044 3000 393096 3052
rect 475108 3000 475160 3052
rect 476948 3000 477000 3052
rect 485688 3000 485740 3052
rect 487620 3000 487672 3052
rect 493968 3000 494020 3052
rect 495900 3000 495952 3052
rect 496912 3000 496964 3052
rect 500592 3000 500644 3052
rect 28908 2932 28960 2984
rect 34888 2932 34940 2984
rect 35992 2932 36044 2984
rect 43352 2932 43404 2984
rect 46664 2932 46716 2984
rect 53104 2932 53156 2984
rect 56048 2932 56100 2984
rect 62672 2932 62724 2984
rect 66720 2932 66772 2984
rect 73160 2932 73212 2984
rect 124680 2932 124732 2984
rect 132408 2932 132460 2984
rect 132960 2932 133012 2984
rect 139584 2932 139636 2984
rect 147128 2932 147180 2984
rect 153200 2932 153252 2984
rect 156604 2932 156656 2984
rect 161480 2932 161532 2984
rect 287244 2932 287296 2984
rect 288992 2932 289044 2984
rect 375380 2932 375432 2984
rect 383568 2932 383620 2984
rect 384396 2932 384448 2984
rect 391848 2932 391900 2984
rect 484676 2932 484728 2984
rect 486424 2932 486476 2984
rect 539692 2932 539744 2984
rect 545488 2932 545540 2984
rect 86868 2864 86920 2916
rect 92480 2864 92532 2916
rect 93952 2864 94004 2916
rect 100944 2864 100996 2916
rect 105728 2864 105780 2916
rect 111984 2864 112036 2916
rect 153016 2864 153068 2916
rect 158720 2864 158772 2916
rect 336740 2864 336792 2916
rect 342168 2864 342220 2916
rect 349068 2864 349120 2916
rect 354036 2864 354088 2916
rect 495348 2864 495400 2916
rect 497096 2864 497148 2916
rect 528652 2864 528704 2916
rect 534908 2864 534960 2916
<< metal2 >>
rect 6932 703582 7972 703610
rect 3422 697368 3478 697377
rect 3422 697303 3478 697312
rect 3436 670682 3464 697303
rect 3514 684312 3570 684321
rect 3514 684247 3570 684256
rect 3424 670676 3476 670682
rect 3424 670618 3476 670624
rect 3528 658238 3556 684247
rect 6932 681018 6960 703582
rect 7944 703474 7972 703582
rect 8086 703520 8198 704960
rect 23492 703582 24164 703610
rect 8128 703474 8156 703520
rect 7944 703446 8156 703474
rect 23492 681018 23520 703582
rect 24136 703474 24164 703582
rect 24278 703520 24390 704960
rect 40052 703582 40356 703610
rect 24320 703474 24348 703520
rect 24136 703446 24348 703474
rect 40052 681018 40080 703582
rect 40328 703474 40356 703582
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218072 703582 218836 703610
rect 40512 703474 40540 703520
rect 40328 703446 40540 703474
rect 56796 683114 56824 703520
rect 72988 703050 73016 703520
rect 71780 703044 71832 703050
rect 71780 702986 71832 702992
rect 72976 703044 73028 703050
rect 72976 702986 73028 702992
rect 56612 683086 56824 683114
rect 56612 681018 56640 683086
rect 71792 681018 71820 702986
rect 89180 702434 89208 703520
rect 88352 702406 89208 702434
rect 88352 681018 88380 702406
rect 105464 699786 105492 703520
rect 105452 699780 105504 699786
rect 105452 699722 105504 699728
rect 108304 699780 108356 699786
rect 108304 699722 108356 699728
rect 6920 681012 6972 681018
rect 6920 680954 6972 680960
rect 19892 681012 19944 681018
rect 19892 680954 19944 680960
rect 23480 681012 23532 681018
rect 23480 680954 23532 680960
rect 35256 681012 35308 681018
rect 35256 680954 35308 680960
rect 40040 681012 40092 681018
rect 40040 680954 40092 680960
rect 50620 681012 50672 681018
rect 50620 680954 50672 680960
rect 56600 681012 56652 681018
rect 56600 680954 56652 680960
rect 66260 681012 66312 681018
rect 66260 680954 66312 680960
rect 71780 681012 71832 681018
rect 71780 680954 71832 680960
rect 81440 681012 81492 681018
rect 81440 680954 81492 680960
rect 88340 681012 88392 681018
rect 88340 680954 88392 680960
rect 96712 681012 96764 681018
rect 96712 680954 96764 680960
rect 19904 678722 19932 680954
rect 35268 678722 35296 680954
rect 50632 678722 50660 680954
rect 66272 678722 66300 680954
rect 81452 678722 81480 680954
rect 96724 678722 96752 680954
rect 108316 680610 108344 699722
rect 121656 699718 121684 703520
rect 137848 699718 137876 703520
rect 154132 699718 154160 703520
rect 170324 699718 170352 703520
rect 186516 699718 186544 703520
rect 202800 699718 202828 703520
rect 121644 699712 121696 699718
rect 121644 699654 121696 699660
rect 124864 699712 124916 699718
rect 124864 699654 124916 699660
rect 137836 699712 137888 699718
rect 137836 699654 137888 699660
rect 140044 699712 140096 699718
rect 140044 699654 140096 699660
rect 154120 699712 154172 699718
rect 154120 699654 154172 699660
rect 156604 699712 156656 699718
rect 156604 699654 156656 699660
rect 170312 699712 170364 699718
rect 170312 699654 170364 699660
rect 172520 699712 172572 699718
rect 172520 699654 172572 699660
rect 186504 699712 186556 699718
rect 186504 699654 186556 699660
rect 189080 699712 189132 699718
rect 189080 699654 189132 699660
rect 202788 699712 202840 699718
rect 202788 699654 202840 699660
rect 204260 699712 204312 699718
rect 204260 699654 204312 699660
rect 108304 680604 108356 680610
rect 108304 680546 108356 680552
rect 112076 680604 112128 680610
rect 112076 680546 112128 680552
rect 112088 678722 112116 680546
rect 124876 680474 124904 699654
rect 140056 680814 140084 699654
rect 140044 680808 140096 680814
rect 140044 680750 140096 680756
rect 142804 680808 142856 680814
rect 142804 680750 142856 680756
rect 124864 680468 124916 680474
rect 124864 680410 124916 680416
rect 127440 680468 127492 680474
rect 127440 680410 127492 680416
rect 127452 678722 127480 680410
rect 142816 678722 142844 680750
rect 156616 680610 156644 699654
rect 172532 692774 172560 699654
rect 172532 692746 173480 692774
rect 156604 680604 156656 680610
rect 156604 680546 156656 680552
rect 158168 680604 158220 680610
rect 158168 680546 158220 680552
rect 158180 678722 158208 680546
rect 173452 678722 173480 692746
rect 189092 678722 189120 699654
rect 204272 678722 204300 699654
rect 218072 680610 218100 703582
rect 218808 703474 218836 703582
rect 218950 703520 219062 704960
rect 234632 703582 235028 703610
rect 218992 703474 219020 703520
rect 218808 703446 219020 703474
rect 234632 692774 234660 703582
rect 235000 703474 235028 703582
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 235184 703474 235212 703520
rect 235000 703446 235212 703474
rect 251468 699718 251496 703520
rect 267660 699718 267688 703520
rect 283852 699718 283880 703520
rect 300136 699718 300164 703520
rect 316328 699718 316356 703520
rect 332520 699718 332548 703520
rect 348804 700330 348832 703520
rect 364996 702434 365024 703520
rect 364352 702406 365024 702434
rect 342260 700324 342312 700330
rect 342260 700266 342312 700272
rect 348792 700324 348844 700330
rect 348792 700266 348844 700272
rect 249800 699712 249852 699718
rect 249800 699654 249852 699660
rect 251456 699712 251508 699718
rect 251456 699654 251508 699660
rect 264980 699712 265032 699718
rect 264980 699654 265032 699660
rect 267648 699712 267700 699718
rect 267648 699654 267700 699660
rect 280160 699712 280212 699718
rect 280160 699654 280212 699660
rect 283840 699712 283892 699718
rect 283840 699654 283892 699660
rect 296720 699712 296772 699718
rect 296720 699654 296772 699660
rect 300124 699712 300176 699718
rect 300124 699654 300176 699660
rect 311900 699712 311952 699718
rect 311900 699654 311952 699660
rect 316316 699712 316368 699718
rect 316316 699654 316368 699660
rect 327080 699712 327132 699718
rect 327080 699654 327132 699660
rect 332508 699712 332560 699718
rect 332508 699654 332560 699660
rect 249812 692774 249840 699654
rect 264992 692774 265020 699654
rect 280172 692774 280200 699654
rect 234632 692746 234936 692774
rect 249812 692746 250300 692774
rect 264992 692746 265664 692774
rect 280172 692746 281028 692774
rect 218060 680604 218112 680610
rect 218060 680546 218112 680552
rect 219716 680604 219768 680610
rect 219716 680546 219768 680552
rect 219728 678722 219756 680546
rect 234908 678722 234936 692746
rect 250272 678722 250300 692746
rect 265636 678722 265664 692746
rect 281000 678722 281028 692746
rect 296732 678722 296760 699654
rect 311912 678722 311940 699654
rect 327092 678722 327120 699654
rect 342272 692774 342300 700266
rect 342272 692746 342484 692774
rect 342456 678722 342484 692746
rect 364352 680746 364380 702406
rect 381188 700330 381216 703520
rect 397472 700330 397500 703520
rect 413664 700330 413692 703520
rect 429856 700330 429884 703520
rect 446140 700330 446168 703520
rect 462332 700330 462360 703520
rect 478524 700330 478552 703520
rect 494808 700330 494836 703520
rect 511000 700466 511028 703520
rect 495440 700460 495492 700466
rect 495440 700402 495492 700408
rect 510988 700460 511040 700466
rect 510988 700402 511040 700408
rect 372620 700324 372672 700330
rect 372620 700266 372672 700272
rect 381176 700324 381228 700330
rect 381176 700266 381228 700272
rect 387800 700324 387852 700330
rect 387800 700266 387852 700272
rect 397460 700324 397512 700330
rect 397460 700266 397512 700272
rect 402980 700324 403032 700330
rect 402980 700266 403032 700272
rect 413652 700324 413704 700330
rect 413652 700266 413704 700272
rect 419540 700324 419592 700330
rect 419540 700266 419592 700272
rect 429844 700324 429896 700330
rect 429844 700266 429896 700272
rect 434720 700324 434772 700330
rect 434720 700266 434772 700272
rect 446128 700324 446180 700330
rect 446128 700266 446180 700272
rect 449900 700324 449952 700330
rect 449900 700266 449952 700272
rect 462320 700324 462372 700330
rect 462320 700266 462372 700272
rect 465080 700324 465132 700330
rect 465080 700266 465132 700272
rect 478512 700324 478564 700330
rect 478512 700266 478564 700272
rect 480260 700324 480312 700330
rect 480260 700266 480312 700272
rect 494796 700324 494848 700330
rect 494796 700266 494848 700272
rect 372632 692774 372660 700266
rect 387812 692774 387840 700266
rect 402992 692774 403020 700266
rect 372632 692746 373212 692774
rect 387812 692746 388576 692774
rect 402992 692746 403940 692774
rect 358544 680740 358596 680746
rect 358544 680682 358596 680688
rect 364340 680740 364392 680746
rect 364340 680682 364392 680688
rect 358556 678722 358584 680682
rect 19904 678694 20240 678722
rect 35268 678694 35604 678722
rect 50632 678694 50968 678722
rect 66272 678694 66332 678722
rect 81452 678694 81696 678722
rect 96724 678694 97060 678722
rect 112088 678694 112424 678722
rect 127452 678694 127788 678722
rect 142816 678694 143152 678722
rect 158180 678694 158516 678722
rect 173452 678694 173880 678722
rect 189092 678694 189244 678722
rect 204272 678694 204608 678722
rect 219728 678694 219972 678722
rect 234908 678694 235336 678722
rect 250272 678694 250700 678722
rect 265636 678694 266064 678722
rect 281000 678694 281428 678722
rect 296732 678694 296792 678722
rect 311912 678694 312156 678722
rect 327092 678694 327520 678722
rect 342456 678694 342884 678722
rect 358248 678694 358584 678722
rect 373184 678722 373212 692746
rect 388548 678722 388576 692746
rect 403912 678722 403940 692746
rect 419552 678722 419580 700266
rect 434732 678722 434760 700266
rect 449912 692774 449940 700266
rect 465092 692774 465120 700266
rect 480272 692774 480300 700266
rect 495452 692774 495480 700402
rect 527192 700330 527220 703520
rect 543476 700534 543504 703520
rect 527272 700528 527324 700534
rect 527272 700470 527324 700476
rect 543464 700528 543516 700534
rect 543464 700470 543516 700476
rect 510620 700324 510672 700330
rect 510620 700266 510672 700272
rect 527180 700324 527232 700330
rect 527180 700266 527232 700272
rect 510632 692774 510660 700266
rect 449912 692746 450032 692774
rect 465092 692746 465396 692774
rect 480272 692746 480760 692774
rect 495452 692746 496124 692774
rect 510632 692746 511488 692774
rect 450004 678722 450032 692746
rect 465368 678722 465396 692746
rect 480732 678722 480760 692746
rect 496096 678722 496124 692746
rect 511460 678722 511488 692746
rect 527284 678994 527312 700470
rect 559668 700398 559696 703520
rect 542360 700392 542412 700398
rect 542360 700334 542412 700340
rect 559656 700392 559708 700398
rect 559656 700334 559708 700340
rect 527238 678966 527312 678994
rect 373184 678694 373612 678722
rect 388548 678694 388976 678722
rect 403912 678694 404340 678722
rect 419552 678694 419704 678722
rect 434732 678694 435068 678722
rect 450004 678694 450432 678722
rect 465368 678694 465796 678722
rect 480732 678694 481160 678722
rect 496096 678694 496524 678722
rect 511460 678694 511888 678722
rect 527238 678708 527266 678966
rect 542372 678722 542400 700334
rect 575860 700330 575888 703520
rect 557540 700324 557592 700330
rect 557540 700266 557592 700272
rect 575848 700324 575900 700330
rect 575848 700266 575900 700272
rect 557552 678722 557580 700266
rect 580170 697232 580226 697241
rect 580170 697167 580226 697176
rect 580184 696998 580212 697167
rect 569224 696992 569276 696998
rect 569224 696934 569276 696940
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 542372 678694 542616 678722
rect 557552 678694 557980 678722
rect 3606 671256 3662 671265
rect 3606 671191 3662 671200
rect 3516 658232 3568 658238
rect 3422 658200 3478 658209
rect 3516 658174 3568 658180
rect 3422 658135 3478 658144
rect 3436 633418 3464 658135
rect 3620 645862 3648 671191
rect 9404 670676 9456 670682
rect 9404 670618 9456 670624
rect 9416 669633 9444 670618
rect 569236 670585 569264 696934
rect 580170 683904 580226 683913
rect 580170 683839 580226 683848
rect 580184 683194 580212 683839
rect 569316 683188 569368 683194
rect 569316 683130 569368 683136
rect 580172 683188 580224 683194
rect 580172 683130 580224 683136
rect 569222 670576 569278 670585
rect 569222 670511 569278 670520
rect 9402 669624 9458 669633
rect 9402 669559 9458 669568
rect 9404 658232 9456 658238
rect 9404 658174 9456 658180
rect 9416 657393 9444 658174
rect 569328 658073 569356 683130
rect 569408 670744 569460 670750
rect 580172 670744 580224 670750
rect 569408 670686 569460 670692
rect 580170 670712 580172 670721
rect 580224 670712 580226 670721
rect 569314 658064 569370 658073
rect 569314 657999 569370 658008
rect 9402 657384 9458 657393
rect 9402 657319 9458 657328
rect 569224 656940 569276 656946
rect 569224 656882 569276 656888
rect 3608 645856 3660 645862
rect 3608 645798 3660 645804
rect 9404 645856 9456 645862
rect 9404 645798 9456 645804
rect 9416 645153 9444 645798
rect 3514 645144 3570 645153
rect 3514 645079 3570 645088
rect 9402 645144 9458 645153
rect 9402 645079 9458 645088
rect 3424 633412 3476 633418
rect 3424 633354 3476 633360
rect 3528 620974 3556 645079
rect 8668 633412 8720 633418
rect 8668 633354 8720 633360
rect 8680 632913 8708 633354
rect 569236 633049 569264 656882
rect 569420 645561 569448 670686
rect 580170 670647 580226 670656
rect 580170 657384 580226 657393
rect 580170 657319 580226 657328
rect 580184 656946 580212 657319
rect 580172 656940 580224 656946
rect 580172 656882 580224 656888
rect 569406 645552 569462 645561
rect 569406 645487 569462 645496
rect 580170 644056 580226 644065
rect 580170 643991 580226 644000
rect 580184 643142 580212 643991
rect 569316 643136 569368 643142
rect 569316 643078 569368 643084
rect 580172 643136 580224 643142
rect 580172 643078 580224 643084
rect 569222 633040 569278 633049
rect 569222 632975 569278 632984
rect 8666 632904 8722 632913
rect 8666 632839 8722 632848
rect 3606 632088 3662 632097
rect 3606 632023 3662 632032
rect 3516 620968 3568 620974
rect 3516 620910 3568 620916
rect 3422 619168 3478 619177
rect 3422 619103 3478 619112
rect 3436 596154 3464 619103
rect 3620 607986 3648 632023
rect 569224 630692 569276 630698
rect 569224 630634 569276 630640
rect 8668 620968 8720 620974
rect 8668 620910 8720 620916
rect 8680 620673 8708 620910
rect 8666 620664 8722 620673
rect 8666 620599 8722 620608
rect 9402 608424 9458 608433
rect 9402 608359 9458 608368
rect 9416 607986 9444 608359
rect 569236 608025 569264 630634
rect 569328 620537 569356 643078
rect 580170 630864 580226 630873
rect 580170 630799 580226 630808
rect 580184 630698 580212 630799
rect 580172 630692 580224 630698
rect 580172 630634 580224 630640
rect 569314 620528 569370 620537
rect 569314 620463 569370 620472
rect 580170 617536 580226 617545
rect 580170 617471 580226 617480
rect 580184 616894 580212 617471
rect 569316 616888 569368 616894
rect 569316 616830 569368 616836
rect 580172 616888 580224 616894
rect 580172 616830 580224 616836
rect 569222 608016 569278 608025
rect 3608 607980 3660 607986
rect 3608 607922 3660 607928
rect 9404 607980 9456 607986
rect 569222 607951 569278 607960
rect 9404 607922 9456 607928
rect 3514 606112 3570 606121
rect 3514 606047 3570 606056
rect 3424 596148 3476 596154
rect 3424 596090 3476 596096
rect 2778 593056 2834 593065
rect 2778 592991 2834 593000
rect 2792 592074 2820 592991
rect 2780 592068 2832 592074
rect 2780 592010 2832 592016
rect 3528 585138 3556 606047
rect 9402 596184 9458 596193
rect 9402 596119 9404 596128
rect 9456 596119 9458 596128
rect 9404 596090 9456 596096
rect 569328 595513 569356 616830
rect 580170 604208 580226 604217
rect 580170 604143 580226 604152
rect 580184 603158 580212 604143
rect 569408 603152 569460 603158
rect 569408 603094 569460 603100
rect 580172 603152 580224 603158
rect 580172 603094 580224 603100
rect 569314 595504 569370 595513
rect 569314 595439 569370 595448
rect 6276 592068 6328 592074
rect 6276 592010 6328 592016
rect 3516 585132 3568 585138
rect 3516 585074 3568 585080
rect 2962 580000 3018 580009
rect 2962 579935 3018 579944
rect 2976 579698 3004 579935
rect 2964 579692 3016 579698
rect 2964 579634 3016 579640
rect 6184 579692 6236 579698
rect 6184 579634 6236 579640
rect 3422 566944 3478 566953
rect 3422 566879 3478 566888
rect 3436 547874 3464 566879
rect 6196 559842 6224 579634
rect 6288 572694 6316 592010
rect 569224 590708 569276 590714
rect 569224 590650 569276 590656
rect 9404 585132 9456 585138
rect 9404 585074 9456 585080
rect 9416 583953 9444 585074
rect 9402 583944 9458 583953
rect 9402 583879 9458 583888
rect 6276 572688 6328 572694
rect 6276 572630 6328 572636
rect 8852 572688 8904 572694
rect 8852 572630 8904 572636
rect 8864 571713 8892 572630
rect 8850 571704 8906 571713
rect 8850 571639 8906 571648
rect 569236 570489 569264 590650
rect 569420 583001 569448 603094
rect 579802 591016 579858 591025
rect 579802 590951 579858 590960
rect 579816 590714 579844 590951
rect 579804 590708 579856 590714
rect 579804 590650 579856 590656
rect 569406 582992 569462 583001
rect 569406 582927 569462 582936
rect 580170 577688 580226 577697
rect 580170 577623 580226 577632
rect 580184 576910 580212 577623
rect 569316 576904 569368 576910
rect 569316 576846 569368 576852
rect 580172 576904 580224 576910
rect 580172 576846 580224 576852
rect 569222 570480 569278 570489
rect 569222 570415 569278 570424
rect 569224 563100 569276 563106
rect 569224 563042 569276 563048
rect 6184 559836 6236 559842
rect 6184 559778 6236 559784
rect 9404 559836 9456 559842
rect 9404 559778 9456 559784
rect 9416 559473 9444 559778
rect 9402 559464 9458 559473
rect 9402 559399 9458 559408
rect 3514 553888 3570 553897
rect 3514 553823 3570 553832
rect 3424 547868 3476 547874
rect 3424 547810 3476 547816
rect 3422 540832 3478 540841
rect 3422 540767 3478 540776
rect 3436 539646 3464 540767
rect 3424 539640 3476 539646
rect 3424 539582 3476 539588
rect 3528 535430 3556 553823
rect 9404 547868 9456 547874
rect 9404 547810 9456 547816
rect 9416 547233 9444 547810
rect 9402 547224 9458 547233
rect 9402 547159 9458 547168
rect 569236 545465 569264 563042
rect 569328 557977 569356 576846
rect 579802 564360 579858 564369
rect 579802 564295 579858 564304
rect 579816 563106 579844 564295
rect 579804 563100 579856 563106
rect 579804 563042 579856 563048
rect 569314 557968 569370 557977
rect 569314 557903 569370 557912
rect 580170 551168 580226 551177
rect 580170 551103 580226 551112
rect 580184 550662 580212 551103
rect 569316 550656 569368 550662
rect 569316 550598 569368 550604
rect 580172 550656 580224 550662
rect 580172 550598 580224 550604
rect 569222 545456 569278 545465
rect 569222 545391 569278 545400
rect 7656 539640 7708 539646
rect 7656 539582 7708 539588
rect 3516 535424 3568 535430
rect 3516 535366 3568 535372
rect 3422 527912 3478 527921
rect 3422 527847 3478 527856
rect 3436 527202 3464 527847
rect 3424 527196 3476 527202
rect 3424 527138 3476 527144
rect 7564 527196 7616 527202
rect 7564 527138 7616 527144
rect 3422 514856 3478 514865
rect 3422 514791 3424 514800
rect 3476 514791 3478 514800
rect 3424 514762 3476 514768
rect 7576 510513 7604 527138
rect 7668 522753 7696 539582
rect 569224 536852 569276 536858
rect 569224 536794 569276 536800
rect 9404 535424 9456 535430
rect 9404 535366 9456 535372
rect 9416 534993 9444 535366
rect 9402 534984 9458 534993
rect 9402 534919 9458 534928
rect 7654 522744 7710 522753
rect 7654 522679 7710 522688
rect 569236 520441 569264 536794
rect 569328 532953 569356 550598
rect 580170 537840 580226 537849
rect 580170 537775 580226 537784
rect 580184 536858 580212 537775
rect 580172 536852 580224 536858
rect 580172 536794 580224 536800
rect 569314 532944 569370 532953
rect 569314 532879 569370 532888
rect 580170 524512 580226 524521
rect 569316 524476 569368 524482
rect 580170 524447 580172 524456
rect 569316 524418 569368 524424
rect 580224 524447 580226 524456
rect 580172 524418 580224 524424
rect 569222 520432 569278 520441
rect 569222 520367 569278 520376
rect 8944 514820 8996 514826
rect 8944 514762 8996 514768
rect 7562 510504 7618 510513
rect 7562 510439 7618 510448
rect 3054 501800 3110 501809
rect 3054 501735 3110 501744
rect 3068 501022 3096 501735
rect 3056 501016 3108 501022
rect 3056 500958 3108 500964
rect 8956 498273 8984 514762
rect 569224 510672 569276 510678
rect 569224 510614 569276 510620
rect 9036 501016 9088 501022
rect 9036 500958 9088 500964
rect 8942 498264 8998 498273
rect 8942 498199 8998 498208
rect 3422 488744 3478 488753
rect 3422 488679 3424 488688
rect 3476 488679 3478 488688
rect 8944 488708 8996 488714
rect 3424 488650 3476 488656
rect 8944 488650 8996 488656
rect 3422 475688 3478 475697
rect 3422 475623 3424 475632
rect 3476 475623 3478 475632
rect 3424 475594 3476 475600
rect 8956 473793 8984 488650
rect 9048 486033 9076 500958
rect 569236 495417 569264 510614
rect 569328 507929 569356 524418
rect 580170 511320 580226 511329
rect 580170 511255 580226 511264
rect 580184 510678 580212 511255
rect 580172 510672 580224 510678
rect 580172 510614 580224 510620
rect 569314 507920 569370 507929
rect 569314 507855 569370 507864
rect 579894 497992 579950 498001
rect 579894 497927 579950 497936
rect 579908 496874 579936 497927
rect 577504 496868 577556 496874
rect 577504 496810 577556 496816
rect 579896 496868 579948 496874
rect 579896 496810 579948 496816
rect 569222 495408 569278 495417
rect 569222 495343 569278 495352
rect 9034 486024 9090 486033
rect 9034 485959 9090 485968
rect 577516 483002 577544 496810
rect 580630 484664 580686 484673
rect 580630 484599 580686 484608
rect 580644 484430 580672 484599
rect 577596 484424 577648 484430
rect 577596 484366 577648 484372
rect 580632 484424 580684 484430
rect 580632 484366 580684 484372
rect 569868 482996 569920 483002
rect 569868 482938 569920 482944
rect 577504 482996 577556 483002
rect 577504 482938 577556 482944
rect 569880 482905 569908 482938
rect 569866 482896 569922 482905
rect 569866 482831 569922 482840
rect 9036 475652 9088 475658
rect 9036 475594 9088 475600
rect 8942 473784 8998 473793
rect 8942 473719 8998 473728
rect 3422 462632 3478 462641
rect 3422 462567 3424 462576
rect 3476 462567 3478 462576
rect 8944 462596 8996 462602
rect 3424 462538 3476 462544
rect 8944 462538 8996 462544
rect 2778 449576 2834 449585
rect 2778 449511 2834 449520
rect 2792 449478 2820 449511
rect 2780 449472 2832 449478
rect 2780 449414 2832 449420
rect 6276 449472 6328 449478
rect 6276 449414 6328 449420
rect 6288 437442 6316 449414
rect 8956 449313 8984 462538
rect 9048 461553 9076 475594
rect 576124 470620 576176 470626
rect 576124 470562 576176 470568
rect 569868 470552 569920 470558
rect 569868 470494 569920 470500
rect 569880 470393 569908 470494
rect 569866 470384 569922 470393
rect 569866 470319 569922 470328
rect 9034 461544 9090 461553
rect 9034 461479 9090 461488
rect 576136 457910 576164 470562
rect 577608 470558 577636 484366
rect 579986 471472 580042 471481
rect 579986 471407 580042 471416
rect 580000 470626 580028 471407
rect 579988 470620 580040 470626
rect 579988 470562 580040 470568
rect 577596 470552 577648 470558
rect 577596 470494 577648 470500
rect 580262 458144 580318 458153
rect 580262 458079 580318 458088
rect 569868 457904 569920 457910
rect 569866 457872 569868 457881
rect 576124 457904 576176 457910
rect 569920 457872 569922 457881
rect 576124 457846 576176 457852
rect 569866 457807 569922 457816
rect 8942 449304 8998 449313
rect 8942 449239 8998 449248
rect 580276 445738 580304 458079
rect 569132 445732 569184 445738
rect 569132 445674 569184 445680
rect 580264 445732 580316 445738
rect 580264 445674 580316 445680
rect 569144 445369 569172 445674
rect 569130 445360 569186 445369
rect 569130 445295 569186 445304
rect 580354 444816 580410 444825
rect 580354 444751 580410 444760
rect 6276 437436 6328 437442
rect 6276 437378 6328 437384
rect 9404 437436 9456 437442
rect 9404 437378 9456 437384
rect 9416 437073 9444 437378
rect 9402 437064 9458 437073
rect 9402 436999 9458 437008
rect 2962 436656 3018 436665
rect 2962 436591 3018 436600
rect 2976 436218 3004 436591
rect 2964 436212 3016 436218
rect 2964 436154 3016 436160
rect 6184 436212 6236 436218
rect 6184 436154 6236 436160
rect 6196 424454 6224 436154
rect 580368 433294 580396 444751
rect 569316 433288 569368 433294
rect 569316 433230 569368 433236
rect 580356 433288 580408 433294
rect 580356 433230 580408 433236
rect 569328 432857 569356 433230
rect 569314 432848 569370 432857
rect 569314 432783 569370 432792
rect 580170 431624 580226 431633
rect 580170 431559 580226 431568
rect 580184 430642 580212 431559
rect 569224 430636 569276 430642
rect 569224 430578 569276 430584
rect 580172 430636 580224 430642
rect 580172 430578 580224 430584
rect 9402 424824 9458 424833
rect 9402 424759 9458 424768
rect 9416 424454 9444 424759
rect 6184 424448 6236 424454
rect 6184 424390 6236 424396
rect 9404 424448 9456 424454
rect 9404 424390 9456 424396
rect 3422 423600 3478 423609
rect 3422 423535 3478 423544
rect 3436 423230 3464 423535
rect 3424 423224 3476 423230
rect 3424 423166 3476 423172
rect 7564 423224 7616 423230
rect 7564 423166 7616 423172
rect 7576 412593 7604 423166
rect 569236 420345 569264 430578
rect 569222 420336 569278 420345
rect 569222 420271 569278 420280
rect 580170 418296 580226 418305
rect 580170 418231 580226 418240
rect 580184 418198 580212 418231
rect 569224 418192 569276 418198
rect 569224 418134 569276 418140
rect 580172 418192 580224 418198
rect 580172 418134 580224 418140
rect 7562 412584 7618 412593
rect 7562 412519 7618 412528
rect 3146 410544 3202 410553
rect 3146 410479 3202 410488
rect 3160 409902 3188 410479
rect 3148 409896 3200 409902
rect 3148 409838 3200 409844
rect 7564 409896 7616 409902
rect 7564 409838 7616 409844
rect 7576 400353 7604 409838
rect 569236 407833 569264 418134
rect 569222 407824 569278 407833
rect 569222 407759 569278 407768
rect 580170 404968 580226 404977
rect 580170 404903 580226 404912
rect 580184 404394 580212 404903
rect 574744 404388 574796 404394
rect 574744 404330 574796 404336
rect 580172 404388 580224 404394
rect 580172 404330 580224 404336
rect 7562 400344 7618 400353
rect 7562 400279 7618 400288
rect 3424 397520 3476 397526
rect 3422 397488 3424 397497
rect 7564 397520 7616 397526
rect 3476 397488 3478 397497
rect 7564 397462 7616 397468
rect 3422 397423 3478 397432
rect 7576 388113 7604 397462
rect 574756 395826 574784 404330
rect 569132 395820 569184 395826
rect 569132 395762 569184 395768
rect 574744 395820 574796 395826
rect 574744 395762 574796 395768
rect 569144 395321 569172 395762
rect 569130 395312 569186 395321
rect 569130 395247 569186 395256
rect 578882 391776 578938 391785
rect 578882 391711 578938 391720
rect 7562 388104 7618 388113
rect 7562 388039 7618 388048
rect 3422 384432 3478 384441
rect 3422 384367 3478 384376
rect 3436 383858 3464 384367
rect 3424 383852 3476 383858
rect 3424 383794 3476 383800
rect 7564 383852 7616 383858
rect 7564 383794 7616 383800
rect 7576 375873 7604 383794
rect 578896 383654 578924 391711
rect 569868 383648 569920 383654
rect 569868 383590 569920 383596
rect 578884 383648 578936 383654
rect 578884 383590 578936 383596
rect 569880 382809 569908 383590
rect 569866 382800 569922 382809
rect 569866 382735 569922 382744
rect 578882 378448 578938 378457
rect 578882 378383 578938 378392
rect 7562 375864 7618 375873
rect 7562 375799 7618 375808
rect 3422 371376 3478 371385
rect 3422 371311 3424 371320
rect 3476 371311 3478 371320
rect 7564 371340 7616 371346
rect 3424 371282 3476 371288
rect 7564 371282 7616 371288
rect 7576 363633 7604 371282
rect 578896 371210 578924 378383
rect 569592 371204 569644 371210
rect 569592 371146 569644 371152
rect 578884 371204 578936 371210
rect 578884 371146 578936 371152
rect 569604 370297 569632 371146
rect 569590 370288 569646 370297
rect 569590 370223 569646 370232
rect 579618 365120 579674 365129
rect 579618 365055 579674 365064
rect 579632 364750 579660 365055
rect 578240 364744 578292 364750
rect 578240 364686 578292 364692
rect 579620 364744 579672 364750
rect 579620 364686 579672 364692
rect 7562 363624 7618 363633
rect 7562 363559 7618 363568
rect 578252 358766 578280 364686
rect 569684 358760 569736 358766
rect 569684 358702 569736 358708
rect 578240 358760 578292 358766
rect 578240 358702 578292 358708
rect 2778 358456 2834 358465
rect 2778 358391 2834 358400
rect 2792 357746 2820 358391
rect 569696 357785 569724 358702
rect 569682 357776 569738 357785
rect 2780 357740 2832 357746
rect 2780 357682 2832 357688
rect 4804 357740 4856 357746
rect 569682 357711 569738 357720
rect 4804 357682 4856 357688
rect 4816 351898 4844 357682
rect 579526 351928 579582 351937
rect 4804 351892 4856 351898
rect 4804 351834 4856 351840
rect 8668 351892 8720 351898
rect 579526 351863 579582 351872
rect 8668 351834 8720 351840
rect 8680 351393 8708 351834
rect 8666 351384 8722 351393
rect 8666 351319 8722 351328
rect 579540 346390 579568 351863
rect 569684 346384 569736 346390
rect 569684 346326 569736 346332
rect 579528 346384 579580 346390
rect 579528 346326 579580 346332
rect 4066 345400 4122 345409
rect 4122 345358 4200 345386
rect 4066 345335 4122 345344
rect 4172 339454 4200 345358
rect 569696 345273 569724 346326
rect 569682 345264 569738 345273
rect 569682 345199 569738 345208
rect 4160 339448 4212 339454
rect 4160 339390 4212 339396
rect 9404 339448 9456 339454
rect 9404 339390 9456 339396
rect 9416 339153 9444 339390
rect 9402 339144 9458 339153
rect 9402 339079 9458 339088
rect 580170 338600 580226 338609
rect 580170 338535 580226 338544
rect 580184 338162 580212 338535
rect 569224 338156 569276 338162
rect 569224 338098 569276 338104
rect 580172 338156 580224 338162
rect 580172 338098 580224 338104
rect 569236 332761 569264 338098
rect 569222 332752 569278 332761
rect 569222 332687 569278 332696
rect 3054 332344 3110 332353
rect 3054 332279 3110 332288
rect 3068 327078 3096 332279
rect 3056 327072 3108 327078
rect 3056 327014 3108 327020
rect 9404 327072 9456 327078
rect 9404 327014 9456 327020
rect 9416 326913 9444 327014
rect 9402 326904 9458 326913
rect 9402 326839 9458 326848
rect 580170 325272 580226 325281
rect 580170 325207 580226 325216
rect 580184 321570 580212 325207
rect 568672 321564 568724 321570
rect 568672 321506 568724 321512
rect 580172 321564 580224 321570
rect 580172 321506 580224 321512
rect 568684 320249 568712 321506
rect 568670 320240 568726 320249
rect 568670 320175 568726 320184
rect 3422 319288 3478 319297
rect 3422 319223 3478 319232
rect 3436 314634 3464 319223
rect 9402 314664 9458 314673
rect 3424 314628 3476 314634
rect 9402 314599 9404 314608
rect 3424 314570 3476 314576
rect 9456 314599 9458 314608
rect 9404 314570 9456 314576
rect 580170 312080 580226 312089
rect 580170 312015 580226 312024
rect 580184 311914 580212 312015
rect 568948 311908 569000 311914
rect 568948 311850 569000 311856
rect 580172 311908 580224 311914
rect 580172 311850 580224 311856
rect 568960 307737 568988 311850
rect 568946 307728 569002 307737
rect 568946 307663 569002 307672
rect 3422 306232 3478 306241
rect 3422 306167 3424 306176
rect 3476 306167 3478 306176
rect 9404 306196 9456 306202
rect 3424 306138 3476 306144
rect 9404 306138 9456 306144
rect 9416 302433 9444 306138
rect 9402 302424 9458 302433
rect 9402 302359 9458 302368
rect 580354 298752 580410 298761
rect 580354 298687 580410 298696
rect 580368 295322 580396 298687
rect 569868 295316 569920 295322
rect 569868 295258 569920 295264
rect 580356 295316 580408 295322
rect 580356 295258 580408 295264
rect 569880 295225 569908 295258
rect 569866 295216 569922 295225
rect 569866 295151 569922 295160
rect 3422 293176 3478 293185
rect 3422 293111 3478 293120
rect 3436 292602 3464 293111
rect 3424 292596 3476 292602
rect 3424 292538 3476 292544
rect 9404 292596 9456 292602
rect 9404 292538 9456 292544
rect 9416 290193 9444 292538
rect 9402 290184 9458 290193
rect 9402 290119 9458 290128
rect 580170 285424 580226 285433
rect 580170 285359 580226 285368
rect 580184 284374 580212 285359
rect 572720 284368 572772 284374
rect 572720 284310 572772 284316
rect 580172 284368 580224 284374
rect 580172 284310 580224 284316
rect 572732 282742 572760 284310
rect 569868 282736 569920 282742
rect 569866 282704 569868 282713
rect 572720 282736 572772 282742
rect 569920 282704 569922 282713
rect 572720 282678 572772 282684
rect 569866 282639 569922 282648
rect 3422 280120 3478 280129
rect 3422 280055 3478 280064
rect 3436 279750 3464 280055
rect 3424 279744 3476 279750
rect 3424 279686 3476 279692
rect 9220 279744 9272 279750
rect 9220 279686 9272 279692
rect 9232 277953 9260 279686
rect 9218 277944 9274 277953
rect 9218 277879 9274 277888
rect 579802 272232 579858 272241
rect 579802 272167 579858 272176
rect 579816 271930 579844 272167
rect 572720 271924 572772 271930
rect 572720 271866 572772 271872
rect 579804 271924 579856 271930
rect 579804 271866 579856 271872
rect 572732 270230 572760 271866
rect 569316 270224 569368 270230
rect 569314 270192 569316 270201
rect 572720 270224 572772 270230
rect 569368 270192 569370 270201
rect 572720 270166 572772 270172
rect 569314 270127 569370 270136
rect 3054 267200 3110 267209
rect 3054 267135 3110 267144
rect 3068 266422 3096 267135
rect 3056 266416 3108 266422
rect 3056 266358 3108 266364
rect 9404 266416 9456 266422
rect 9404 266358 9456 266364
rect 9416 265713 9444 266358
rect 9402 265704 9458 265713
rect 9402 265639 9458 265648
rect 579710 258904 579766 258913
rect 579710 258839 579766 258848
rect 579724 258126 579752 258839
rect 579712 258120 579764 258126
rect 579712 258062 579764 258068
rect 569132 258052 569184 258058
rect 569132 257994 569184 258000
rect 569144 257689 569172 257994
rect 569130 257680 569186 257689
rect 569130 257615 569186 257624
rect 3422 254144 3478 254153
rect 3422 254079 3424 254088
rect 3476 254079 3478 254088
rect 9404 254108 9456 254114
rect 3424 254050 3476 254056
rect 9404 254050 9456 254056
rect 9416 253473 9444 254050
rect 9402 253464 9458 253473
rect 9402 253399 9458 253408
rect 580170 245576 580226 245585
rect 580170 245511 580226 245520
rect 568670 245168 568726 245177
rect 568670 245103 568726 245112
rect 568684 244934 568712 245103
rect 580184 244934 580212 245511
rect 568672 244928 568724 244934
rect 568672 244870 568724 244876
rect 580172 244928 580224 244934
rect 580172 244870 580224 244876
rect 9402 241224 9458 241233
rect 9402 241159 9458 241168
rect 3422 241088 3478 241097
rect 3422 241023 3478 241032
rect 3436 240922 3464 241023
rect 9416 240922 9444 241159
rect 3424 240916 3476 240922
rect 3424 240858 3476 240864
rect 9404 240916 9456 240922
rect 9404 240858 9456 240864
rect 569866 232656 569922 232665
rect 569866 232591 569922 232600
rect 569880 232558 569908 232591
rect 569868 232552 569920 232558
rect 569868 232494 569920 232500
rect 580172 232552 580224 232558
rect 580172 232494 580224 232500
rect 580184 232393 580212 232494
rect 580170 232384 580226 232393
rect 580170 232319 580226 232328
rect 8850 228984 8906 228993
rect 8850 228919 8906 228928
rect 3422 228032 3478 228041
rect 8864 228002 8892 228919
rect 3422 227967 3424 227976
rect 3476 227967 3478 227976
rect 8852 227996 8904 228002
rect 3424 227938 3476 227944
rect 8852 227938 8904 227944
rect 569498 220144 569554 220153
rect 569498 220079 569554 220088
rect 569512 219502 569540 220079
rect 569500 219496 569552 219502
rect 569500 219438 569552 219444
rect 580448 219428 580500 219434
rect 580448 219370 580500 219376
rect 580460 219065 580488 219370
rect 580446 219056 580502 219065
rect 580446 218991 580502 219000
rect 8206 216744 8262 216753
rect 8206 216679 8262 216688
rect 8220 215014 8248 216679
rect 3424 215008 3476 215014
rect 3422 214976 3424 214985
rect 8208 215008 8260 215014
rect 3476 214976 3478 214985
rect 8208 214950 8260 214956
rect 3422 214911 3478 214920
rect 569866 207632 569922 207641
rect 569866 207567 569922 207576
rect 569880 207058 569908 207567
rect 569868 207052 569920 207058
rect 569868 206994 569920 207000
rect 579528 207052 579580 207058
rect 579528 206994 579580 207000
rect 579540 205737 579568 206994
rect 579526 205728 579582 205737
rect 579526 205663 579582 205672
rect 8206 204504 8262 204513
rect 8206 204439 8262 204448
rect 8220 202230 8248 204439
rect 3332 202224 3384 202230
rect 3332 202166 3384 202172
rect 8208 202224 8260 202230
rect 8208 202166 8260 202172
rect 3344 201929 3372 202166
rect 3330 201920 3386 201929
rect 3330 201855 3386 201864
rect 569314 195120 569370 195129
rect 569314 195055 569370 195064
rect 569328 194614 569356 195055
rect 569316 194608 569368 194614
rect 569316 194550 569368 194556
rect 579528 194608 579580 194614
rect 579528 194550 579580 194556
rect 579540 192545 579568 194550
rect 579526 192536 579582 192545
rect 579526 192471 579582 192480
rect 8206 192264 8262 192273
rect 8206 192199 8262 192208
rect 8220 188902 8248 192199
rect 3424 188896 3476 188902
rect 3422 188864 3424 188873
rect 8208 188896 8260 188902
rect 3476 188864 3478 188873
rect 8208 188838 8260 188844
rect 3422 188799 3478 188808
rect 569406 182608 569462 182617
rect 569406 182543 569462 182552
rect 569420 182238 569448 182543
rect 569408 182232 569460 182238
rect 569408 182174 569460 182180
rect 576860 182232 576912 182238
rect 576860 182174 576912 182180
rect 8206 180024 8262 180033
rect 8206 179959 8262 179968
rect 8220 176662 8248 179959
rect 576872 179382 576900 182174
rect 576860 179376 576912 179382
rect 576860 179318 576912 179324
rect 580264 179376 580316 179382
rect 580264 179318 580316 179324
rect 580276 179217 580304 179318
rect 580262 179208 580318 179217
rect 580262 179143 580318 179152
rect 3424 176656 3476 176662
rect 3424 176598 3476 176604
rect 8208 176656 8260 176662
rect 8208 176598 8260 176604
rect 3436 175953 3464 176598
rect 3422 175944 3478 175953
rect 3422 175879 3478 175888
rect 569866 170096 569922 170105
rect 569866 170031 569922 170040
rect 569880 169794 569908 170031
rect 569868 169788 569920 169794
rect 569868 169730 569920 169736
rect 577964 169788 578016 169794
rect 577964 169730 578016 169736
rect 8206 167784 8262 167793
rect 8206 167719 8262 167728
rect 8220 163402 8248 167719
rect 577976 167006 578004 169730
rect 577964 167000 578016 167006
rect 577964 166942 578016 166948
rect 579988 167000 580040 167006
rect 579988 166942 580040 166948
rect 580000 165889 580028 166942
rect 579986 165880 580042 165889
rect 579986 165815 580042 165824
rect 3516 163396 3568 163402
rect 3516 163338 3568 163344
rect 8208 163396 8260 163402
rect 8208 163338 8260 163344
rect 3528 162897 3556 163338
rect 3514 162888 3570 162897
rect 3514 162823 3570 162832
rect 569866 157584 569922 157593
rect 569866 157519 569922 157528
rect 569880 157418 569908 157519
rect 569868 157412 569920 157418
rect 569868 157354 569920 157360
rect 579528 157412 579580 157418
rect 579528 157354 579580 157360
rect 8942 155544 8998 155553
rect 8942 155479 8998 155488
rect 8956 150414 8984 155479
rect 579540 152697 579568 157354
rect 579526 152688 579582 152697
rect 579526 152623 579582 152632
rect 3424 150408 3476 150414
rect 3424 150350 3476 150356
rect 8944 150408 8996 150414
rect 8944 150350 8996 150356
rect 3436 149841 3464 150350
rect 3422 149832 3478 149841
rect 3422 149767 3478 149776
rect 569866 145072 569922 145081
rect 569866 145007 569922 145016
rect 569880 144974 569908 145007
rect 569868 144968 569920 144974
rect 569868 144910 569920 144916
rect 578884 144968 578936 144974
rect 578884 144910 578936 144916
rect 8298 143304 8354 143313
rect 8298 143239 8354 143248
rect 8312 137970 8340 143239
rect 578896 139369 578924 144910
rect 578882 139360 578938 139369
rect 578882 139295 578938 139304
rect 3240 137964 3292 137970
rect 3240 137906 3292 137912
rect 8300 137964 8352 137970
rect 8300 137906 8352 137912
rect 3252 136785 3280 137906
rect 3238 136776 3294 136785
rect 3238 136711 3294 136720
rect 569866 132560 569922 132569
rect 569866 132495 569868 132504
rect 569920 132495 569922 132504
rect 578240 132524 578292 132530
rect 569868 132466 569920 132472
rect 578240 132466 578292 132472
rect 9034 131064 9090 131073
rect 9034 130999 9090 131008
rect 9048 129810 9076 130999
rect 4160 129804 4212 129810
rect 4160 129746 4212 129752
rect 9036 129804 9088 129810
rect 9036 129746 9088 129752
rect 4066 123720 4122 123729
rect 4172 123706 4200 129746
rect 578252 126954 578280 132466
rect 578240 126948 578292 126954
rect 578240 126890 578292 126896
rect 579620 126948 579672 126954
rect 579620 126890 579672 126896
rect 579632 126041 579660 126890
rect 579618 126032 579674 126041
rect 579618 125967 579674 125976
rect 4122 123678 4200 123706
rect 4066 123655 4122 123664
rect 568670 120048 568726 120057
rect 568670 119983 568726 119992
rect 9402 118824 9458 118833
rect 9402 118759 9458 118768
rect 9416 118726 9444 118759
rect 568684 118726 568712 119983
rect 4804 118720 4856 118726
rect 4804 118662 4856 118668
rect 9404 118720 9456 118726
rect 9404 118662 9456 118668
rect 568672 118720 568724 118726
rect 568672 118662 568724 118668
rect 578884 118720 578936 118726
rect 578884 118662 578936 118668
rect 4816 110770 4844 118662
rect 578896 112849 578924 118662
rect 578882 112840 578938 112849
rect 578882 112775 578938 112784
rect 2780 110764 2832 110770
rect 2780 110706 2832 110712
rect 4804 110764 4856 110770
rect 4804 110706 4856 110712
rect 2792 110673 2820 110706
rect 2778 110664 2834 110673
rect 2778 110599 2834 110608
rect 569682 107536 569738 107545
rect 569682 107471 569738 107480
rect 9402 106584 9458 106593
rect 9402 106519 9458 106528
rect 9416 106350 9444 106519
rect 569696 106350 569724 107471
rect 4804 106344 4856 106350
rect 4804 106286 4856 106292
rect 9404 106344 9456 106350
rect 9404 106286 9456 106292
rect 569684 106344 569736 106350
rect 569684 106286 569736 106292
rect 578884 106344 578936 106350
rect 578884 106286 578936 106292
rect 4816 97782 4844 106286
rect 578896 99521 578924 106286
rect 578882 99512 578938 99521
rect 578882 99447 578938 99456
rect 2780 97776 2832 97782
rect 2780 97718 2832 97724
rect 4804 97776 4856 97782
rect 4804 97718 4856 97724
rect 2792 97617 2820 97718
rect 2778 97608 2834 97617
rect 2778 97543 2834 97552
rect 569682 95024 569738 95033
rect 569682 94959 569738 94968
rect 569696 94450 569724 94959
rect 569684 94444 569736 94450
rect 569684 94386 569736 94392
rect 576124 94444 576176 94450
rect 576124 94386 576176 94392
rect 9402 94344 9458 94353
rect 9402 94279 9458 94288
rect 9416 93906 9444 94279
rect 4804 93900 4856 93906
rect 4804 93842 4856 93848
rect 9404 93900 9456 93906
rect 9404 93842 9456 93848
rect 4816 85270 4844 93842
rect 576136 86970 576164 94386
rect 576124 86964 576176 86970
rect 576124 86906 576176 86912
rect 580172 86964 580224 86970
rect 580172 86906 580224 86912
rect 580184 86193 580212 86906
rect 580170 86184 580226 86193
rect 580170 86119 580226 86128
rect 2780 85264 2832 85270
rect 2780 85206 2832 85212
rect 4804 85264 4856 85270
rect 4804 85206 4856 85212
rect 2792 84697 2820 85206
rect 2778 84688 2834 84697
rect 2778 84623 2834 84632
rect 569682 82512 569738 82521
rect 569682 82447 569738 82456
rect 8942 82104 8998 82113
rect 8942 82039 8998 82048
rect 8956 71670 8984 82039
rect 569696 81462 569724 82447
rect 569684 81456 569736 81462
rect 569684 81398 569736 81404
rect 578884 81456 578936 81462
rect 578884 81398 578936 81404
rect 578896 73001 578924 81398
rect 578882 72992 578938 73001
rect 578882 72927 578938 72936
rect 3424 71664 3476 71670
rect 3422 71632 3424 71641
rect 8944 71664 8996 71670
rect 3476 71632 3478 71641
rect 8944 71606 8996 71612
rect 3422 71567 3478 71576
rect 569590 70000 569646 70009
rect 569590 69935 569646 69944
rect 8942 69864 8998 69873
rect 8942 69799 8998 69808
rect 8956 59226 8984 69799
rect 569604 69086 569632 69935
rect 569592 69080 569644 69086
rect 569592 69022 569644 69028
rect 578884 69080 578936 69086
rect 578884 69022 578936 69028
rect 578896 59673 578924 69022
rect 578882 59664 578938 59673
rect 578882 59599 578938 59608
rect 3148 59220 3200 59226
rect 3148 59162 3200 59168
rect 8944 59220 8996 59226
rect 8944 59162 8996 59168
rect 3160 58585 3188 59162
rect 3146 58576 3202 58585
rect 3146 58511 3202 58520
rect 8850 57624 8906 57633
rect 8850 57559 8906 57568
rect 8864 56642 8892 57559
rect 569130 57488 569186 57497
rect 569130 57423 569186 57432
rect 569144 56642 569172 57423
rect 4804 56636 4856 56642
rect 4804 56578 4856 56584
rect 8852 56636 8904 56642
rect 8852 56578 8904 56584
rect 569132 56636 569184 56642
rect 569132 56578 569184 56584
rect 574744 56636 574796 56642
rect 574744 56578 574796 56584
rect 4816 45558 4844 56578
rect 574756 46918 574784 56578
rect 574744 46912 574796 46918
rect 574744 46854 574796 46860
rect 580172 46912 580224 46918
rect 580172 46854 580224 46860
rect 580184 46345 580212 46854
rect 580170 46336 580226 46345
rect 580170 46271 580226 46280
rect 2780 45552 2832 45558
rect 2778 45520 2780 45529
rect 4804 45552 4856 45558
rect 2832 45520 2834 45529
rect 4804 45494 4856 45500
rect 2778 45455 2834 45464
rect 9402 45384 9458 45393
rect 9402 45319 9458 45328
rect 9416 44198 9444 45319
rect 569866 44976 569922 44985
rect 569866 44911 569922 44920
rect 569880 44198 569908 44911
rect 4896 44192 4948 44198
rect 4896 44134 4948 44140
rect 9404 44192 9456 44198
rect 9404 44134 9456 44140
rect 569868 44192 569920 44198
rect 569868 44134 569920 44140
rect 578884 44192 578936 44198
rect 578884 44134 578936 44140
rect 4908 32910 4936 44134
rect 578896 33153 578924 44134
rect 9034 33144 9090 33153
rect 9034 33079 9090 33088
rect 578882 33144 578938 33153
rect 578882 33079 578938 33088
rect 2780 32904 2832 32910
rect 2780 32846 2832 32852
rect 4896 32904 4948 32910
rect 4896 32846 4948 32852
rect 2792 32473 2820 32846
rect 2778 32464 2834 32473
rect 2778 32399 2834 32408
rect 9048 31822 9076 33079
rect 569498 32464 569554 32473
rect 569498 32399 569554 32408
rect 569512 31822 569540 32399
rect 4804 31816 4856 31822
rect 4804 31758 4856 31764
rect 9036 31816 9088 31822
rect 9036 31758 9088 31764
rect 569500 31816 569552 31822
rect 569500 31758 569552 31764
rect 578976 31816 579028 31822
rect 578976 31758 579028 31764
rect 4816 20398 4844 31758
rect 8942 20904 8998 20913
rect 8942 20839 8998 20848
rect 2780 20392 2832 20398
rect 2780 20334 2832 20340
rect 4804 20392 4856 20398
rect 4804 20334 4856 20340
rect 2792 19417 2820 20334
rect 2778 19408 2834 19417
rect 2778 19343 2834 19352
rect 8956 6526 8984 20839
rect 569866 19952 569922 19961
rect 569866 19887 569922 19896
rect 569880 19378 569908 19887
rect 578988 19825 579016 31758
rect 578974 19816 579030 19825
rect 578974 19751 579030 19760
rect 569868 19372 569920 19378
rect 569868 19314 569920 19320
rect 578884 19372 578936 19378
rect 578884 19314 578936 19320
rect 16684 12022 16928 12050
rect 18032 12022 18184 12050
rect 15200 8968 15252 8974
rect 15200 8910 15252 8916
rect 13820 8356 13872 8362
rect 13820 8298 13872 8304
rect 3424 6520 3476 6526
rect 3422 6488 3424 6497
rect 8944 6520 8996 6526
rect 3476 6488 3478 6497
rect 8944 6462 8996 6468
rect 3422 6423 3478 6432
rect 5264 4140 5316 4146
rect 5264 4082 5316 4088
rect 4068 3936 4120 3942
rect 4068 3878 4120 3884
rect 2872 3868 2924 3874
rect 2872 3810 2924 3816
rect 572 3800 624 3806
rect 572 3742 624 3748
rect 584 480 612 3742
rect 1676 3460 1728 3466
rect 1676 3402 1728 3408
rect 1688 480 1716 3402
rect 2884 480 2912 3810
rect 4080 480 4108 3878
rect 5276 480 5304 4082
rect 9956 4004 10008 4010
rect 9956 3946 10008 3952
rect 6460 3664 6512 3670
rect 6460 3606 6512 3612
rect 6472 480 6500 3606
rect 7656 3528 7708 3534
rect 7656 3470 7708 3476
rect 7668 480 7696 3470
rect 8760 3324 8812 3330
rect 8760 3266 8812 3272
rect 8772 480 8800 3266
rect 9968 480 9996 3946
rect 13832 3806 13860 8298
rect 15212 4146 15240 8910
rect 16684 8362 16712 12022
rect 17960 9512 18012 9518
rect 17960 9454 18012 9460
rect 17868 9172 17920 9178
rect 17868 9114 17920 9120
rect 16672 8356 16724 8362
rect 16672 8298 16724 8304
rect 16764 8356 16816 8362
rect 16764 8298 16816 8304
rect 16776 6914 16804 8298
rect 16684 6886 16804 6914
rect 15200 4140 15252 4146
rect 15200 4082 15252 4088
rect 14740 4072 14792 4078
rect 14740 4014 14792 4020
rect 13820 3800 13872 3806
rect 13820 3742 13872 3748
rect 11152 3732 11204 3738
rect 11152 3674 11204 3680
rect 11164 480 11192 3674
rect 12348 3596 12400 3602
rect 12348 3538 12400 3544
rect 12360 480 12388 3538
rect 13544 3392 13596 3398
rect 13544 3334 13596 3340
rect 13556 480 13584 3334
rect 14752 480 14780 4014
rect 16684 3942 16712 6886
rect 16672 3936 16724 3942
rect 16672 3878 16724 3884
rect 17880 3874 17908 9114
rect 17868 3868 17920 3874
rect 17868 3810 17920 3816
rect 15936 3800 15988 3806
rect 15936 3742 15988 3748
rect 15948 480 15976 3742
rect 17972 3330 18000 9454
rect 18052 3936 18104 3942
rect 18052 3878 18104 3884
rect 18064 3534 18092 3878
rect 18052 3528 18104 3534
rect 18052 3470 18104 3476
rect 18156 3466 18184 12022
rect 18800 12022 19136 12050
rect 19904 12022 20240 12050
rect 21008 12022 21344 12050
rect 22204 12022 22448 12050
rect 23552 12022 23704 12050
rect 18800 9178 18828 12022
rect 18788 9172 18840 9178
rect 18788 9114 18840 9120
rect 19904 8362 19932 12022
rect 21008 8974 21036 12022
rect 20996 8968 21048 8974
rect 20996 8910 21048 8916
rect 22100 8900 22152 8906
rect 22100 8842 22152 8848
rect 19892 8356 19944 8362
rect 19892 8298 19944 8304
rect 22112 4010 22140 8842
rect 22100 4004 22152 4010
rect 22100 3946 22152 3952
rect 21824 3868 21876 3874
rect 21824 3810 21876 3816
rect 18236 3528 18288 3534
rect 18236 3470 18288 3476
rect 18144 3460 18196 3466
rect 18144 3402 18196 3408
rect 17960 3324 18012 3330
rect 17960 3266 18012 3272
rect 17040 3188 17092 3194
rect 17040 3130 17092 3136
rect 17052 480 17080 3130
rect 18248 480 18276 3470
rect 19432 3460 19484 3466
rect 19432 3402 19484 3408
rect 19444 480 19472 3402
rect 20628 3324 20680 3330
rect 20628 3266 20680 3272
rect 20640 480 20668 3266
rect 21836 480 21864 3810
rect 22204 3670 22232 12022
rect 23296 9308 23348 9314
rect 23296 9250 23348 9256
rect 22192 3664 22244 3670
rect 22192 3606 22244 3612
rect 23020 3664 23072 3670
rect 23020 3606 23072 3612
rect 23032 480 23060 3606
rect 23308 3398 23336 9250
rect 23388 9104 23440 9110
rect 23388 9046 23440 9052
rect 23400 3806 23428 9046
rect 23676 3942 23704 12022
rect 24320 12022 24656 12050
rect 25424 12022 25760 12050
rect 26252 12022 26864 12050
rect 27816 12022 27968 12050
rect 29012 12022 29072 12050
rect 29840 12022 30176 12050
rect 30944 12022 31280 12050
rect 32048 12022 32384 12050
rect 33152 12022 33488 12050
rect 34532 12022 34592 12050
rect 35360 12022 35696 12050
rect 36464 12022 36800 12050
rect 37568 12022 37904 12050
rect 38672 12022 39008 12050
rect 40052 12022 40112 12050
rect 40880 12022 41216 12050
rect 41984 12022 42320 12050
rect 43088 12022 43424 12050
rect 44192 12022 44528 12050
rect 45572 12022 45632 12050
rect 46400 12022 46736 12050
rect 47504 12022 47840 12050
rect 48608 12022 48944 12050
rect 49712 12022 50048 12050
rect 51092 12022 51152 12050
rect 51920 12022 52256 12050
rect 53024 12022 53360 12050
rect 54128 12022 54464 12050
rect 55324 12022 55568 12050
rect 56612 12022 56672 12050
rect 57440 12022 57776 12050
rect 58544 12022 58880 12050
rect 59648 12022 59984 12050
rect 60752 12022 61088 12050
rect 62132 12022 62192 12050
rect 62960 12022 63296 12050
rect 64064 12022 64400 12050
rect 65168 12022 65504 12050
rect 66272 12022 66608 12050
rect 67652 12022 67712 12050
rect 68480 12022 68816 12050
rect 69584 12022 69920 12050
rect 70688 12022 71024 12050
rect 71792 12022 72128 12050
rect 73172 12022 73232 12050
rect 74000 12022 74336 12050
rect 75104 12022 75440 12050
rect 76208 12022 76544 12050
rect 77312 12022 77648 12050
rect 78692 12022 78752 12050
rect 79520 12022 79856 12050
rect 80624 12022 80960 12050
rect 81728 12022 82064 12050
rect 82832 12022 83168 12050
rect 84212 12022 84272 12050
rect 85040 12022 85376 12050
rect 86144 12022 86480 12050
rect 87248 12022 87584 12050
rect 88352 12022 88688 12050
rect 89732 12022 89792 12050
rect 90560 12022 90896 12050
rect 91664 12022 92000 12050
rect 92768 12022 93104 12050
rect 93964 12022 94208 12050
rect 95252 12022 95312 12050
rect 96080 12022 96416 12050
rect 97184 12022 97520 12050
rect 98288 12022 98624 12050
rect 99392 12022 99728 12050
rect 100772 12022 100832 12050
rect 101600 12022 101936 12050
rect 102704 12022 103040 12050
rect 103808 12022 104144 12050
rect 104912 12022 105248 12050
rect 106292 12022 106352 12050
rect 107120 12022 107456 12050
rect 108224 12022 108560 12050
rect 109328 12022 109664 12050
rect 110432 12022 110768 12050
rect 111812 12022 111872 12050
rect 112640 12022 112976 12050
rect 113744 12022 114080 12050
rect 114848 12022 115184 12050
rect 115952 12022 116288 12050
rect 117332 12022 117392 12050
rect 118160 12022 118496 12050
rect 119264 12022 119600 12050
rect 120368 12022 120704 12050
rect 121472 12022 121808 12050
rect 24320 9518 24348 12022
rect 24308 9512 24360 9518
rect 24308 9454 24360 9460
rect 24952 9444 25004 9450
rect 24952 9386 25004 9392
rect 24032 9172 24084 9178
rect 24032 9114 24084 9120
rect 23664 3936 23716 3942
rect 23664 3878 23716 3884
rect 23388 3800 23440 3806
rect 23388 3742 23440 3748
rect 23296 3392 23348 3398
rect 23296 3334 23348 3340
rect 24044 3194 24072 9114
rect 24964 4078 24992 9386
rect 25044 9240 25096 9246
rect 25044 9182 25096 9188
rect 24952 4072 25004 4078
rect 24952 4014 25004 4020
rect 24216 4004 24268 4010
rect 24216 3946 24268 3952
rect 24032 3188 24084 3194
rect 24032 3130 24084 3136
rect 24228 480 24256 3946
rect 25056 3534 25084 9182
rect 25424 8906 25452 12022
rect 25412 8900 25464 8906
rect 25412 8842 25464 8848
rect 25320 3800 25372 3806
rect 25320 3742 25372 3748
rect 25044 3528 25096 3534
rect 25044 3470 25096 3476
rect 25332 480 25360 3742
rect 26252 3738 26280 12022
rect 26332 9580 26384 9586
rect 26332 9522 26384 9528
rect 26240 3732 26292 3738
rect 26240 3674 26292 3680
rect 26344 3330 26372 9522
rect 26424 9512 26476 9518
rect 26424 9454 26476 9460
rect 26436 3466 26464 9454
rect 27620 8968 27672 8974
rect 27620 8910 27672 8916
rect 27632 3874 27660 8910
rect 27620 3868 27672 3874
rect 27620 3810 27672 3816
rect 27816 3602 27844 12022
rect 29012 9314 29040 12022
rect 29840 9450 29868 12022
rect 29828 9444 29880 9450
rect 29828 9386 29880 9392
rect 29000 9308 29052 9314
rect 29000 9250 29052 9256
rect 29920 9308 29972 9314
rect 29920 9250 29972 9256
rect 29932 3670 29960 9250
rect 30944 9110 30972 12022
rect 32048 9178 32076 12022
rect 33152 9246 33180 12022
rect 34532 9518 34560 12022
rect 35360 9586 35388 12022
rect 35348 9580 35400 9586
rect 35348 9522 35400 9528
rect 35992 9580 36044 9586
rect 35992 9522 36044 9528
rect 34520 9512 34572 9518
rect 34520 9454 34572 9460
rect 34704 9512 34756 9518
rect 34704 9454 34756 9460
rect 33784 9444 33836 9450
rect 33784 9386 33836 9392
rect 33140 9240 33192 9246
rect 33140 9182 33192 9188
rect 32036 9172 32088 9178
rect 32036 9114 32088 9120
rect 32772 9172 32824 9178
rect 32772 9114 32824 9120
rect 30932 9104 30984 9110
rect 30932 9046 30984 9052
rect 31668 9104 31720 9110
rect 31668 9046 31720 9052
rect 30104 4140 30156 4146
rect 30104 4082 30156 4088
rect 29920 3664 29972 3670
rect 29920 3606 29972 3612
rect 27804 3596 27856 3602
rect 27804 3538 27856 3544
rect 26516 3528 26568 3534
rect 26516 3470 26568 3476
rect 26424 3460 26476 3466
rect 26424 3402 26476 3408
rect 26332 3324 26384 3330
rect 26332 3266 26384 3272
rect 26528 480 26556 3470
rect 27712 3392 27764 3398
rect 27712 3334 27764 3340
rect 27724 480 27752 3334
rect 28908 2984 28960 2990
rect 28908 2926 28960 2932
rect 28920 480 28948 2926
rect 30116 480 30144 4082
rect 31680 4010 31708 9046
rect 31668 4004 31720 4010
rect 31668 3946 31720 3952
rect 31300 3868 31352 3874
rect 31300 3810 31352 3816
rect 31312 480 31340 3810
rect 32784 3806 32812 9114
rect 32772 3800 32824 3806
rect 32772 3742 32824 3748
rect 32404 3732 32456 3738
rect 32404 3674 32456 3680
rect 32416 480 32444 3674
rect 33600 3596 33652 3602
rect 33600 3538 33652 3544
rect 33612 480 33640 3538
rect 33796 3534 33824 9386
rect 33784 3528 33836 3534
rect 33784 3470 33836 3476
rect 34716 3398 34744 9454
rect 34888 9376 34940 9382
rect 34888 9318 34940 9324
rect 34796 3800 34848 3806
rect 34796 3742 34848 3748
rect 34704 3392 34756 3398
rect 34704 3334 34756 3340
rect 34808 480 34836 3742
rect 34900 2990 34928 9318
rect 36004 4146 36032 9522
rect 36464 8974 36492 12022
rect 37568 9314 37596 12022
rect 37556 9308 37608 9314
rect 37556 9250 37608 9256
rect 38672 9110 38700 12022
rect 40052 9178 40080 12022
rect 40880 9450 40908 12022
rect 41984 9518 42012 12022
rect 41972 9512 42024 9518
rect 41972 9454 42024 9460
rect 40868 9444 40920 9450
rect 40868 9386 40920 9392
rect 41328 9444 41380 9450
rect 41328 9386 41380 9392
rect 40040 9172 40092 9178
rect 40040 9114 40092 9120
rect 38660 9104 38712 9110
rect 38660 9046 38712 9052
rect 37280 9036 37332 9042
rect 37280 8978 37332 8984
rect 36452 8968 36504 8974
rect 36452 8910 36504 8916
rect 35992 4140 36044 4146
rect 35992 4082 36044 4088
rect 37292 3874 37320 8978
rect 39304 8356 39356 8362
rect 39304 8298 39356 8304
rect 37280 3868 37332 3874
rect 37280 3810 37332 3816
rect 39316 3738 39344 8298
rect 39580 4140 39632 4146
rect 39580 4082 39632 4088
rect 39304 3732 39356 3738
rect 39304 3674 39356 3680
rect 37188 3528 37240 3534
rect 37188 3470 37240 3476
rect 34888 2984 34940 2990
rect 34888 2926 34940 2932
rect 35992 2984 36044 2990
rect 35992 2926 36044 2932
rect 36004 480 36032 2926
rect 37200 480 37228 3470
rect 38384 3052 38436 3058
rect 38384 2994 38436 3000
rect 38396 480 38424 2994
rect 39592 480 39620 4082
rect 41340 3602 41368 9386
rect 43088 9382 43116 12022
rect 44192 9586 44220 12022
rect 44180 9580 44232 9586
rect 44180 9522 44232 9528
rect 43076 9376 43128 9382
rect 43076 9318 43128 9324
rect 43352 9376 43404 9382
rect 43352 9318 43404 9324
rect 41512 9172 41564 9178
rect 41512 9114 41564 9120
rect 41524 3806 41552 9114
rect 41512 3800 41564 3806
rect 41512 3742 41564 3748
rect 43076 3800 43128 3806
rect 43076 3742 43128 3748
rect 41880 3732 41932 3738
rect 41880 3674 41932 3680
rect 41328 3596 41380 3602
rect 41328 3538 41380 3544
rect 40684 3324 40736 3330
rect 40684 3266 40736 3272
rect 40696 480 40724 3266
rect 41892 480 41920 3674
rect 43088 480 43116 3742
rect 43364 2990 43392 9318
rect 44364 9240 44416 9246
rect 44364 9182 44416 9188
rect 43444 8968 43496 8974
rect 43444 8910 43496 8916
rect 43456 3534 43484 8910
rect 44272 3936 44324 3942
rect 44272 3878 44324 3884
rect 43444 3528 43496 3534
rect 43444 3470 43496 3476
rect 43352 2984 43404 2990
rect 43352 2926 43404 2932
rect 44284 480 44312 3878
rect 44376 3058 44404 9182
rect 45572 9042 45600 12022
rect 45744 9512 45796 9518
rect 45744 9454 45796 9460
rect 45560 9036 45612 9042
rect 45560 8978 45612 8984
rect 45756 4146 45784 9454
rect 46400 8362 46428 12022
rect 47504 9450 47532 12022
rect 47492 9444 47544 9450
rect 47492 9386 47544 9392
rect 46940 9308 46992 9314
rect 46940 9250 46992 9256
rect 46388 8356 46440 8362
rect 46388 8298 46440 8304
rect 45744 4140 45796 4146
rect 45744 4082 45796 4088
rect 45468 3460 45520 3466
rect 45468 3402 45520 3408
rect 44364 3052 44416 3058
rect 44364 2994 44416 3000
rect 45480 480 45508 3402
rect 46952 3330 46980 9250
rect 48608 9178 48636 12022
rect 49712 9382 49740 12022
rect 49700 9376 49752 9382
rect 49700 9318 49752 9324
rect 50988 9376 51040 9382
rect 50988 9318 51040 9324
rect 48596 9172 48648 9178
rect 48596 9114 48648 9120
rect 49608 9172 49660 9178
rect 49608 9114 49660 9120
rect 49620 3738 49648 9114
rect 50160 4140 50212 4146
rect 50160 4082 50212 4088
rect 49608 3732 49660 3738
rect 49608 3674 49660 3680
rect 47860 3528 47912 3534
rect 47860 3470 47912 3476
rect 46940 3324 46992 3330
rect 46940 3266 46992 3272
rect 46664 2984 46716 2990
rect 46664 2926 46716 2932
rect 46676 480 46704 2926
rect 47872 480 47900 3470
rect 48964 3324 49016 3330
rect 48964 3266 49016 3272
rect 48976 480 49004 3266
rect 50172 480 50200 4082
rect 51000 3806 51028 9318
rect 51092 8974 51120 12022
rect 51920 9246 51948 12022
rect 53024 9518 53052 12022
rect 53012 9512 53064 9518
rect 53012 9454 53064 9460
rect 52276 9444 52328 9450
rect 52276 9386 52328 9392
rect 51908 9240 51960 9246
rect 51908 9182 51960 9188
rect 51080 8968 51132 8974
rect 51080 8910 51132 8916
rect 52092 8356 52144 8362
rect 52092 8298 52144 8304
rect 52104 3942 52132 8298
rect 52092 3936 52144 3942
rect 52092 3878 52144 3884
rect 50988 3800 51040 3806
rect 50988 3742 51040 3748
rect 51356 3800 51408 3806
rect 51356 3742 51408 3748
rect 51368 480 51396 3742
rect 52288 3466 52316 9386
rect 54128 9314 54156 12022
rect 54116 9308 54168 9314
rect 54116 9250 54168 9256
rect 53932 9240 53984 9246
rect 53932 9182 53984 9188
rect 53104 8968 53156 8974
rect 53104 8910 53156 8916
rect 52276 3460 52328 3466
rect 52276 3402 52328 3408
rect 52552 3460 52604 3466
rect 52552 3402 52604 3408
rect 52564 480 52592 3402
rect 53116 2990 53144 8910
rect 53748 4072 53800 4078
rect 53748 4014 53800 4020
rect 53104 2984 53156 2990
rect 53104 2926 53156 2932
rect 53760 480 53788 4014
rect 53944 3534 53972 9182
rect 55324 9178 55352 12022
rect 56612 9382 56640 12022
rect 56600 9376 56652 9382
rect 56600 9318 56652 9324
rect 56692 9308 56744 9314
rect 56692 9250 56744 9256
rect 55312 9172 55364 9178
rect 55312 9114 55364 9120
rect 55220 8900 55272 8906
rect 55220 8842 55272 8848
rect 54944 4004 54996 4010
rect 54944 3946 54996 3952
rect 53932 3528 53984 3534
rect 53932 3470 53984 3476
rect 54956 480 54984 3946
rect 55232 3330 55260 8842
rect 56704 4146 56732 9250
rect 57440 8362 57468 12022
rect 58544 9450 58572 12022
rect 58532 9444 58584 9450
rect 58532 9386 58584 9392
rect 59268 9444 59320 9450
rect 59268 9386 59320 9392
rect 57428 8356 57480 8362
rect 57428 8298 57480 8304
rect 56692 4140 56744 4146
rect 56692 4082 56744 4088
rect 58440 4140 58492 4146
rect 58440 4082 58492 4088
rect 57244 3528 57296 3534
rect 57244 3470 57296 3476
rect 55220 3324 55272 3330
rect 55220 3266 55272 3272
rect 56048 2984 56100 2990
rect 56048 2926 56100 2932
rect 56060 480 56088 2926
rect 57256 480 57284 3470
rect 58452 480 58480 4082
rect 59280 3806 59308 9386
rect 59648 8974 59676 12022
rect 60752 9246 60780 12022
rect 60740 9240 60792 9246
rect 60740 9182 60792 9188
rect 59636 8968 59688 8974
rect 59636 8910 59688 8916
rect 60924 8968 60976 8974
rect 60924 8910 60976 8916
rect 60556 8424 60608 8430
rect 60556 8366 60608 8372
rect 60004 8356 60056 8362
rect 60004 8298 60056 8304
rect 60016 4078 60044 8298
rect 60004 4072 60056 4078
rect 60004 4014 60056 4020
rect 59268 3800 59320 3806
rect 59268 3742 59320 3748
rect 59636 3596 59688 3602
rect 59636 3538 59688 3544
rect 59648 480 59676 3538
rect 60568 3466 60596 8366
rect 60936 4010 60964 8910
rect 62132 8906 62160 12022
rect 62960 9314 62988 12022
rect 64064 9450 64092 12022
rect 64052 9444 64104 9450
rect 64052 9386 64104 9392
rect 64972 9376 65024 9382
rect 64972 9318 65024 9324
rect 62948 9308 63000 9314
rect 62948 9250 63000 9256
rect 63500 9308 63552 9314
rect 63500 9250 63552 9256
rect 62672 9172 62724 9178
rect 62672 9114 62724 9120
rect 62120 8900 62172 8906
rect 62120 8842 62172 8848
rect 62028 4072 62080 4078
rect 62028 4014 62080 4020
rect 60924 4004 60976 4010
rect 60924 3946 60976 3952
rect 60556 3460 60608 3466
rect 60556 3402 60608 3408
rect 60832 3460 60884 3466
rect 60832 3402 60884 3408
rect 60844 480 60872 3402
rect 62040 480 62068 4014
rect 62684 2990 62712 9114
rect 63224 3664 63276 3670
rect 63224 3606 63276 3612
rect 62672 2984 62724 2990
rect 62672 2926 62724 2932
rect 63236 480 63264 3606
rect 63512 3534 63540 9250
rect 64984 4146 65012 9318
rect 65168 8430 65196 12022
rect 65156 8424 65208 8430
rect 65156 8366 65208 8372
rect 66272 8362 66300 12022
rect 66352 9444 66404 9450
rect 66352 9386 66404 9392
rect 66260 8356 66312 8362
rect 66260 8298 66312 8304
rect 64972 4140 65024 4146
rect 64972 4082 65024 4088
rect 64328 3800 64380 3806
rect 64328 3742 64380 3748
rect 63500 3528 63552 3534
rect 63500 3470 63552 3476
rect 64340 480 64368 3742
rect 66364 3602 66392 9386
rect 67652 8974 67680 12022
rect 68480 9178 68508 12022
rect 68652 9580 68704 9586
rect 68652 9522 68704 9528
rect 68468 9172 68520 9178
rect 68468 9114 68520 9120
rect 67640 8968 67692 8974
rect 67640 8910 67692 8916
rect 67916 4140 67968 4146
rect 67916 4082 67968 4088
rect 66352 3596 66404 3602
rect 66352 3538 66404 3544
rect 65524 3392 65576 3398
rect 65524 3334 65576 3340
rect 65536 480 65564 3334
rect 66720 2984 66772 2990
rect 66720 2926 66772 2932
rect 66732 480 66760 2926
rect 67928 480 67956 4082
rect 68664 4078 68692 9522
rect 68928 9512 68980 9518
rect 68928 9454 68980 9460
rect 68652 4072 68704 4078
rect 68652 4014 68704 4020
rect 68940 3466 68968 9454
rect 69584 9314 69612 12022
rect 70688 9382 70716 12022
rect 71792 9450 71820 12022
rect 73172 9518 73200 12022
rect 74000 9586 74028 12022
rect 73988 9580 74040 9586
rect 73988 9522 74040 9528
rect 73160 9512 73212 9518
rect 73160 9454 73212 9460
rect 71780 9444 71832 9450
rect 71780 9386 71832 9392
rect 74632 9444 74684 9450
rect 74632 9386 74684 9392
rect 70676 9376 70728 9382
rect 70676 9318 70728 9324
rect 69572 9308 69624 9314
rect 69572 9250 69624 9256
rect 70952 9308 71004 9314
rect 70952 9250 71004 9256
rect 69940 8424 69992 8430
rect 69940 8366 69992 8372
rect 69112 4072 69164 4078
rect 69112 4014 69164 4020
rect 68928 3460 68980 3466
rect 68928 3402 68980 3408
rect 69124 480 69152 4014
rect 69952 3670 69980 8366
rect 70964 3806 70992 9250
rect 72424 9240 72476 9246
rect 72424 9182 72476 9188
rect 71504 3868 71556 3874
rect 71504 3810 71556 3816
rect 70952 3800 71004 3806
rect 70952 3742 71004 3748
rect 69940 3664 69992 3670
rect 69940 3606 69992 3612
rect 70308 3460 70360 3466
rect 70308 3402 70360 3408
rect 70320 480 70348 3402
rect 71516 480 71544 3810
rect 72436 3398 72464 9182
rect 73160 9036 73212 9042
rect 73160 8978 73212 8984
rect 72608 3664 72660 3670
rect 72608 3606 72660 3612
rect 72424 3392 72476 3398
rect 72424 3334 72476 3340
rect 72620 480 72648 3606
rect 73172 2990 73200 8978
rect 74644 4146 74672 9386
rect 75104 8430 75132 12022
rect 75920 9648 75972 9654
rect 75920 9590 75972 9596
rect 75092 8424 75144 8430
rect 75092 8366 75144 8372
rect 74632 4140 74684 4146
rect 74632 4082 74684 4088
rect 73804 3732 73856 3738
rect 73804 3674 73856 3680
rect 73160 2984 73212 2990
rect 73160 2926 73212 2932
rect 73816 480 73844 3674
rect 75000 3528 75052 3534
rect 75000 3470 75052 3476
rect 75012 480 75040 3470
rect 75932 3466 75960 9590
rect 76104 9512 76156 9518
rect 76104 9454 76156 9460
rect 76116 4078 76144 9454
rect 76208 9314 76236 12022
rect 76196 9308 76248 9314
rect 76196 9250 76248 9256
rect 77312 9246 77340 12022
rect 78588 9580 78640 9586
rect 78588 9522 78640 9528
rect 77300 9240 77352 9246
rect 77300 9182 77352 9188
rect 76104 4072 76156 4078
rect 76104 4014 76156 4020
rect 77392 4072 77444 4078
rect 77392 4014 77444 4020
rect 75920 3460 75972 3466
rect 75920 3402 75972 3408
rect 76196 3052 76248 3058
rect 76196 2994 76248 3000
rect 76208 480 76236 2994
rect 77404 480 77432 4014
rect 78600 3874 78628 9522
rect 78692 9042 78720 12022
rect 79520 9450 79548 12022
rect 80624 9518 80652 12022
rect 81728 9654 81756 12022
rect 81716 9648 81768 9654
rect 81716 9590 81768 9596
rect 82832 9586 82860 12022
rect 82820 9580 82872 9586
rect 82820 9522 82872 9528
rect 80612 9512 80664 9518
rect 80612 9454 80664 9460
rect 79508 9444 79560 9450
rect 79508 9386 79560 9392
rect 81532 9376 81584 9382
rect 81532 9318 81584 9324
rect 79968 9308 80020 9314
rect 79968 9250 80020 9256
rect 78680 9036 78732 9042
rect 78680 8978 78732 8984
rect 79692 4140 79744 4146
rect 79692 4082 79744 4088
rect 78588 3868 78640 3874
rect 78588 3810 78640 3816
rect 78588 3324 78640 3330
rect 78588 3266 78640 3272
rect 78600 480 78628 3266
rect 79704 480 79732 4082
rect 79980 3670 80008 9250
rect 80520 8356 80572 8362
rect 80520 8298 80572 8304
rect 80532 3738 80560 8298
rect 80888 3868 80940 3874
rect 80888 3810 80940 3816
rect 80520 3732 80572 3738
rect 80520 3674 80572 3680
rect 79968 3664 80020 3670
rect 79968 3606 80020 3612
rect 80900 480 80928 3810
rect 81544 3534 81572 9318
rect 84212 9314 84240 12022
rect 84384 9512 84436 9518
rect 84384 9454 84436 9460
rect 84200 9308 84252 9314
rect 84200 9250 84252 9256
rect 82820 9104 82872 9110
rect 82820 9046 82872 9052
rect 82084 3596 82136 3602
rect 82084 3538 82136 3544
rect 81532 3528 81584 3534
rect 81532 3470 81584 3476
rect 82096 480 82124 3538
rect 82832 3058 82860 9046
rect 84292 8628 84344 8634
rect 84292 8570 84344 8576
rect 83280 3528 83332 3534
rect 83280 3470 83332 3476
rect 82820 3052 82872 3058
rect 82820 2994 82872 3000
rect 83292 480 83320 3470
rect 84304 3330 84332 8570
rect 84396 4078 84424 9454
rect 85040 8362 85068 12022
rect 86144 9382 86172 12022
rect 86132 9376 86184 9382
rect 86132 9318 86184 9324
rect 87248 9110 87276 12022
rect 88352 9518 88380 12022
rect 88340 9512 88392 9518
rect 88340 9454 88392 9460
rect 89628 9444 89680 9450
rect 89628 9386 89680 9392
rect 87788 9172 87840 9178
rect 87788 9114 87840 9120
rect 87236 9104 87288 9110
rect 87236 9046 87288 9052
rect 85580 8900 85632 8906
rect 85580 8842 85632 8848
rect 85028 8356 85080 8362
rect 85028 8298 85080 8304
rect 85592 4146 85620 8842
rect 85580 4140 85632 4146
rect 85580 4082 85632 4088
rect 84384 4072 84436 4078
rect 84384 4014 84436 4020
rect 87800 3874 87828 9114
rect 89168 4140 89220 4146
rect 89168 4082 89220 4088
rect 87788 3868 87840 3874
rect 87788 3810 87840 3816
rect 85672 3460 85724 3466
rect 85672 3402 85724 3408
rect 84292 3324 84344 3330
rect 84292 3266 84344 3272
rect 84476 3052 84528 3058
rect 84476 2994 84528 3000
rect 84488 480 84516 2994
rect 85684 480 85712 3402
rect 87972 3324 88024 3330
rect 87972 3266 88024 3272
rect 86868 2916 86920 2922
rect 86868 2858 86920 2864
rect 86880 480 86908 2858
rect 87984 480 88012 3266
rect 89180 480 89208 4082
rect 89640 3602 89668 9386
rect 89732 8634 89760 12022
rect 90180 9104 90232 9110
rect 90180 9046 90232 9052
rect 89720 8628 89772 8634
rect 89720 8570 89772 8576
rect 89628 3596 89680 3602
rect 89628 3538 89680 3544
rect 90192 3534 90220 9046
rect 90560 8906 90588 12022
rect 91664 9178 91692 12022
rect 92768 9450 92796 12022
rect 93860 9512 93912 9518
rect 93860 9454 93912 9460
rect 92756 9444 92808 9450
rect 92756 9386 92808 9392
rect 92572 9240 92624 9246
rect 92572 9182 92624 9188
rect 91652 9172 91704 9178
rect 91652 9114 91704 9120
rect 92480 9172 92532 9178
rect 92480 9114 92532 9120
rect 90548 8900 90600 8906
rect 90548 8842 90600 8848
rect 91192 8356 91244 8362
rect 91192 8298 91244 8304
rect 90364 3596 90416 3602
rect 90364 3538 90416 3544
rect 90180 3528 90232 3534
rect 90180 3470 90232 3476
rect 90376 480 90404 3538
rect 91204 3058 91232 8298
rect 91560 3528 91612 3534
rect 91560 3470 91612 3476
rect 91192 3052 91244 3058
rect 91192 2994 91244 3000
rect 91572 480 91600 3470
rect 92492 2922 92520 9114
rect 92584 3466 92612 9182
rect 92756 3732 92808 3738
rect 92756 3674 92808 3680
rect 92572 3460 92624 3466
rect 92572 3402 92624 3408
rect 92480 2916 92532 2922
rect 92480 2858 92532 2864
rect 92768 480 92796 3674
rect 93872 3330 93900 9454
rect 93964 9110 93992 12022
rect 93952 9104 94004 9110
rect 93952 9046 94004 9052
rect 95252 8362 95280 12022
rect 95332 9376 95384 9382
rect 95332 9318 95384 9324
rect 95240 8356 95292 8362
rect 95240 8298 95292 8304
rect 95344 6914 95372 9318
rect 96080 9246 96108 12022
rect 96068 9240 96120 9246
rect 96068 9182 96120 9188
rect 97184 9178 97212 12022
rect 98288 9518 98316 12022
rect 98276 9512 98328 9518
rect 98276 9454 98328 9460
rect 98460 9512 98512 9518
rect 98460 9454 98512 9460
rect 97172 9172 97224 9178
rect 97172 9114 97224 9120
rect 97172 9036 97224 9042
rect 97172 8978 97224 8984
rect 95252 6886 95372 6914
rect 95252 4146 95280 6886
rect 95240 4140 95292 4146
rect 95240 4082 95292 4088
rect 97184 3602 97212 8978
rect 97448 4140 97500 4146
rect 97448 4082 97500 4088
rect 97172 3596 97224 3602
rect 97172 3538 97224 3544
rect 95148 3460 95200 3466
rect 95148 3402 95200 3408
rect 93860 3324 93912 3330
rect 93860 3266 93912 3272
rect 93952 2916 94004 2922
rect 93952 2858 94004 2864
rect 93964 480 93992 2858
rect 95160 480 95188 3402
rect 96252 3392 96304 3398
rect 96252 3334 96304 3340
rect 96264 480 96292 3334
rect 97460 480 97488 4082
rect 98472 3534 98500 9454
rect 99392 9382 99420 12022
rect 99472 9444 99524 9450
rect 99472 9386 99524 9392
rect 99380 9376 99432 9382
rect 99380 9318 99432 9324
rect 99484 3738 99512 9386
rect 100772 9042 100800 12022
rect 101600 9518 101628 12022
rect 101588 9512 101640 9518
rect 101588 9454 101640 9460
rect 102704 9450 102732 12022
rect 103612 9580 103664 9586
rect 103612 9522 103664 9528
rect 102692 9444 102744 9450
rect 102692 9386 102744 9392
rect 100760 9036 100812 9042
rect 100760 8978 100812 8984
rect 102140 9036 102192 9042
rect 102140 8978 102192 8984
rect 100944 8424 100996 8430
rect 100944 8366 100996 8372
rect 100852 8356 100904 8362
rect 100852 8298 100904 8304
rect 99840 3800 99892 3806
rect 99840 3742 99892 3748
rect 99472 3732 99524 3738
rect 99472 3674 99524 3680
rect 98460 3528 98512 3534
rect 98460 3470 98512 3476
rect 98644 3188 98696 3194
rect 98644 3130 98696 3136
rect 98656 480 98684 3130
rect 99852 480 99880 3742
rect 100864 3466 100892 8298
rect 100852 3460 100904 3466
rect 100852 3402 100904 3408
rect 100956 2922 100984 8366
rect 101036 3936 101088 3942
rect 101036 3878 101088 3884
rect 100944 2916 100996 2922
rect 100944 2858 100996 2864
rect 101048 480 101076 3878
rect 102152 3398 102180 8978
rect 103624 4146 103652 9522
rect 103808 8430 103836 12022
rect 103796 8424 103848 8430
rect 103796 8366 103848 8372
rect 104912 8362 104940 12022
rect 104992 9512 105044 9518
rect 104992 9454 105044 9460
rect 104900 8356 104952 8362
rect 104900 8298 104952 8304
rect 103612 4140 103664 4146
rect 103612 4082 103664 4088
rect 104532 3664 104584 3670
rect 104532 3606 104584 3612
rect 103336 3528 103388 3534
rect 103336 3470 103388 3476
rect 102232 3460 102284 3466
rect 102232 3402 102284 3408
rect 102140 3392 102192 3398
rect 102140 3334 102192 3340
rect 102244 480 102272 3402
rect 103348 480 103376 3470
rect 104544 480 104572 3606
rect 105004 3194 105032 9454
rect 106292 9042 106320 12022
rect 107120 9586 107148 12022
rect 107108 9580 107160 9586
rect 107108 9522 107160 9528
rect 108224 9518 108252 12022
rect 109132 9580 109184 9586
rect 109132 9522 109184 9528
rect 108212 9512 108264 9518
rect 108212 9454 108264 9460
rect 106832 9444 106884 9450
rect 106832 9386 106884 9392
rect 106280 9036 106332 9042
rect 106280 8978 106332 8984
rect 106844 3806 106872 9386
rect 108212 8764 108264 8770
rect 108212 8706 108264 8712
rect 108120 4140 108172 4146
rect 108120 4082 108172 4088
rect 106832 3800 106884 3806
rect 106832 3742 106884 3748
rect 106924 3732 106976 3738
rect 106924 3674 106976 3680
rect 104992 3188 105044 3194
rect 104992 3130 105044 3136
rect 105728 2916 105780 2922
rect 105728 2858 105780 2864
rect 105740 480 105768 2858
rect 106936 480 106964 3674
rect 108132 480 108160 4082
rect 108224 3942 108252 8706
rect 108212 3936 108264 3942
rect 108212 3878 108264 3884
rect 109144 3534 109172 9522
rect 109224 9512 109276 9518
rect 109224 9454 109276 9460
rect 109132 3528 109184 3534
rect 109132 3470 109184 3476
rect 109236 3466 109264 9454
rect 109328 9450 109356 12022
rect 109316 9444 109368 9450
rect 109316 9386 109368 9392
rect 110432 8770 110460 12022
rect 111812 9518 111840 12022
rect 112640 9586 112668 12022
rect 112628 9580 112680 9586
rect 112628 9522 112680 9528
rect 111800 9512 111852 9518
rect 111800 9454 111852 9460
rect 113272 9444 113324 9450
rect 113272 9386 113324 9392
rect 111984 9172 112036 9178
rect 111984 9114 112036 9120
rect 110420 8764 110472 8770
rect 110420 8706 110472 8712
rect 110512 8356 110564 8362
rect 110512 8298 110564 8304
rect 110524 3670 110552 8298
rect 111616 4004 111668 4010
rect 111616 3946 111668 3952
rect 110512 3664 110564 3670
rect 110512 3606 110564 3612
rect 109316 3596 109368 3602
rect 109316 3538 109368 3544
rect 109224 3460 109276 3466
rect 109224 3402 109276 3408
rect 109328 480 109356 3538
rect 110512 3460 110564 3466
rect 110512 3402 110564 3408
rect 110524 480 110552 3402
rect 111628 480 111656 3946
rect 111996 2922 112024 9114
rect 113284 3738 113312 9386
rect 113744 8362 113772 12022
rect 114560 9512 114612 9518
rect 114560 9454 114612 9460
rect 113732 8356 113784 8362
rect 113732 8298 113784 8304
rect 114572 4146 114600 9454
rect 114848 9178 114876 12022
rect 115952 9450 115980 12022
rect 117332 9518 117360 12022
rect 117320 9512 117372 9518
rect 117320 9454 117372 9460
rect 118160 9450 118188 12022
rect 119264 9518 119292 12022
rect 118608 9512 118660 9518
rect 118608 9454 118660 9460
rect 119252 9512 119304 9518
rect 119252 9454 119304 9460
rect 115940 9444 115992 9450
rect 115940 9386 115992 9392
rect 117228 9444 117280 9450
rect 117228 9386 117280 9392
rect 118148 9444 118200 9450
rect 118148 9386 118200 9392
rect 114836 9172 114888 9178
rect 114836 9114 114888 9120
rect 114560 4140 114612 4146
rect 114560 4082 114612 4088
rect 116400 4140 116452 4146
rect 116400 4082 116452 4088
rect 113272 3732 113324 3738
rect 113272 3674 113324 3680
rect 112812 3528 112864 3534
rect 112812 3470 112864 3476
rect 111984 2916 112036 2922
rect 111984 2858 112036 2864
rect 112824 480 112852 3470
rect 115204 3392 115256 3398
rect 115204 3334 115256 3340
rect 114008 3052 114060 3058
rect 114008 2994 114060 3000
rect 114020 480 114048 2994
rect 115216 480 115244 3334
rect 116412 480 116440 4082
rect 117240 3602 117268 9386
rect 118056 9036 118108 9042
rect 118056 8978 118108 8984
rect 118068 4010 118096 8978
rect 118056 4004 118108 4010
rect 118056 3946 118108 3952
rect 117228 3596 117280 3602
rect 117228 3538 117280 3544
rect 118620 3466 118648 9454
rect 118700 9444 118752 9450
rect 118700 9386 118752 9392
rect 118712 3534 118740 9386
rect 120368 9042 120396 12022
rect 121472 9450 121500 12022
rect 122898 11778 122926 12036
rect 123680 12022 124016 12050
rect 124784 12022 125120 12050
rect 125888 12022 126224 12050
rect 126992 12022 127328 12050
rect 128372 12022 128432 12050
rect 129200 12022 129536 12050
rect 130304 12022 130640 12050
rect 131132 12022 131744 12050
rect 132512 12022 132848 12050
rect 133892 12022 133952 12050
rect 134168 12022 135056 12050
rect 135824 12022 136160 12050
rect 136652 12022 137264 12050
rect 138032 12022 138368 12050
rect 139412 12022 139472 12050
rect 139596 12022 140576 12050
rect 140792 12022 141680 12050
rect 142172 12022 142784 12050
rect 143552 12022 143888 12050
rect 144932 12022 144992 12050
rect 145116 12022 146096 12050
rect 146312 12022 147200 12050
rect 147692 12022 148304 12050
rect 149072 12022 149408 12050
rect 150452 12022 150512 12050
rect 150636 12022 151616 12050
rect 151832 12022 152720 12050
rect 153212 12022 153824 12050
rect 154592 12022 154928 12050
rect 122898 11750 122972 11778
rect 122760 9654 122880 9674
rect 122760 9648 122892 9654
rect 122760 9646 122840 9648
rect 121460 9444 121512 9450
rect 121460 9386 121512 9392
rect 120356 9036 120408 9042
rect 120356 8978 120408 8984
rect 120172 8356 120224 8362
rect 120172 8298 120224 8304
rect 118792 4004 118844 4010
rect 118792 3946 118844 3952
rect 118700 3528 118752 3534
rect 118700 3470 118752 3476
rect 118608 3460 118660 3466
rect 118608 3402 118660 3408
rect 117596 3324 117648 3330
rect 117596 3266 117648 3272
rect 117608 480 117636 3266
rect 118804 480 118832 3946
rect 119896 3460 119948 3466
rect 119896 3402 119948 3408
rect 119908 480 119936 3402
rect 120184 3058 120212 8298
rect 122288 3868 122340 3874
rect 122288 3810 122340 3816
rect 121092 3732 121144 3738
rect 121092 3674 121144 3680
rect 120172 3052 120224 3058
rect 120172 2994 120224 3000
rect 121104 480 121132 3674
rect 122300 480 122328 3810
rect 122760 3398 122788 9646
rect 122840 9590 122892 9596
rect 122944 8362 122972 11750
rect 123680 9654 123708 12022
rect 123668 9648 123720 9654
rect 123668 9590 123720 9596
rect 124220 9580 124272 9586
rect 124220 9522 124272 9528
rect 124128 9512 124180 9518
rect 124128 9454 124180 9460
rect 122932 8356 122984 8362
rect 122932 8298 122984 8304
rect 124140 4146 124168 9454
rect 124128 4140 124180 4146
rect 124128 4082 124180 4088
rect 122748 3392 122800 3398
rect 122748 3334 122800 3340
rect 124232 3330 124260 9522
rect 124784 9518 124812 12022
rect 125888 9586 125916 12022
rect 125876 9580 125928 9586
rect 125876 9522 125928 9528
rect 124772 9512 124824 9518
rect 124772 9454 124824 9460
rect 126520 8900 126572 8906
rect 126520 8842 126572 8848
rect 125876 4072 125928 4078
rect 125876 4014 125928 4020
rect 124220 3324 124272 3330
rect 124220 3266 124272 3272
rect 123484 3052 123536 3058
rect 123484 2994 123536 3000
rect 123496 480 123524 2994
rect 124680 2984 124732 2990
rect 124680 2926 124732 2932
rect 124692 480 124720 2926
rect 125888 480 125916 4014
rect 126532 3466 126560 8842
rect 126992 8378 127020 12022
rect 128268 9444 128320 9450
rect 128268 9386 128320 9392
rect 126900 8350 127020 8378
rect 126900 4010 126928 8350
rect 128176 4140 128228 4146
rect 128176 4082 128228 4088
rect 126888 4004 126940 4010
rect 126888 3946 126940 3952
rect 126520 3460 126572 3466
rect 126520 3402 126572 3408
rect 126980 3188 127032 3194
rect 126980 3130 127032 3136
rect 126992 480 127020 3130
rect 128188 480 128216 4082
rect 128280 3738 128308 9386
rect 128372 8906 128400 12022
rect 129200 9450 129228 12022
rect 130304 9518 130332 12022
rect 129648 9512 129700 9518
rect 129648 9454 129700 9460
rect 130292 9512 130344 9518
rect 131132 9466 131160 12022
rect 132512 9674 132540 12022
rect 130292 9454 130344 9460
rect 129188 9444 129240 9450
rect 129188 9386 129240 9392
rect 128360 8900 128412 8906
rect 128360 8842 128412 8848
rect 129660 3874 129688 9454
rect 131040 9438 131160 9466
rect 132420 9646 132540 9674
rect 129648 3868 129700 3874
rect 129648 3810 129700 3816
rect 128268 3732 128320 3738
rect 128268 3674 128320 3680
rect 130568 3664 130620 3670
rect 130568 3606 130620 3612
rect 129372 3460 129424 3466
rect 129372 3402 129424 3408
rect 129384 480 129412 3402
rect 130580 480 130608 3606
rect 131040 3058 131068 9438
rect 131764 3596 131816 3602
rect 131764 3538 131816 3544
rect 131028 3052 131080 3058
rect 131028 2994 131080 3000
rect 131776 480 131804 3538
rect 132420 2990 132448 9646
rect 133892 9466 133920 12022
rect 133800 9438 133920 9466
rect 133800 4078 133828 9438
rect 133880 9376 133932 9382
rect 133880 9318 133932 9324
rect 133892 4146 133920 9318
rect 134168 6914 134196 12022
rect 135824 9382 135852 12022
rect 136652 9466 136680 12022
rect 136560 9438 136680 9466
rect 135812 9376 135864 9382
rect 135812 9318 135864 9324
rect 133984 6886 134196 6914
rect 133880 4140 133932 4146
rect 133880 4082 133932 4088
rect 133788 4072 133840 4078
rect 133788 4014 133840 4020
rect 133984 3194 134012 6886
rect 136456 4072 136508 4078
rect 136456 4014 136508 4020
rect 135260 3256 135312 3262
rect 135260 3198 135312 3204
rect 133972 3188 134024 3194
rect 133972 3130 134024 3136
rect 134156 3052 134208 3058
rect 134156 2994 134208 3000
rect 132408 2984 132460 2990
rect 132408 2926 132460 2932
rect 132960 2984 133012 2990
rect 132960 2926 133012 2932
rect 132972 480 133000 2926
rect 134168 480 134196 2994
rect 135272 480 135300 3198
rect 136468 480 136496 4014
rect 136560 3466 136588 9438
rect 138032 8378 138060 12022
rect 139412 9466 139440 12022
rect 137940 8350 138060 8378
rect 139320 9438 139440 9466
rect 137652 4140 137704 4146
rect 137652 4082 137704 4088
rect 136548 3460 136600 3466
rect 136548 3402 136600 3408
rect 137664 480 137692 4082
rect 137940 3670 137968 8350
rect 137928 3664 137980 3670
rect 137928 3606 137980 3612
rect 138848 3664 138900 3670
rect 138848 3606 138900 3612
rect 138860 480 138888 3606
rect 139320 3602 139348 9438
rect 139308 3596 139360 3602
rect 139308 3538 139360 3544
rect 139596 2990 139624 12022
rect 140044 3732 140096 3738
rect 140044 3674 140096 3680
rect 139584 2984 139636 2990
rect 139584 2926 139636 2932
rect 140056 480 140084 3674
rect 140792 3058 140820 12022
rect 141240 3868 141292 3874
rect 141240 3810 141292 3816
rect 140780 3052 140832 3058
rect 140780 2994 140832 3000
rect 141252 480 141280 3810
rect 142172 3262 142200 12022
rect 143552 9466 143580 12022
rect 143460 9438 143580 9466
rect 143460 4078 143488 9438
rect 144932 9382 144960 12022
rect 143540 9376 143592 9382
rect 143540 9318 143592 9324
rect 144920 9376 144972 9382
rect 144920 9318 144972 9324
rect 143552 4146 143580 9318
rect 143540 4140 143592 4146
rect 143540 4082 143592 4088
rect 143448 4072 143500 4078
rect 143448 4014 143500 4020
rect 145116 3670 145144 12022
rect 145932 4140 145984 4146
rect 145932 4082 145984 4088
rect 145104 3664 145156 3670
rect 145104 3606 145156 3612
rect 142436 3460 142488 3466
rect 142436 3402 142488 3408
rect 142160 3256 142212 3262
rect 142160 3198 142212 3204
rect 142448 480 142476 3402
rect 143540 3324 143592 3330
rect 143540 3266 143592 3272
rect 143552 480 143580 3266
rect 144736 3052 144788 3058
rect 144736 2994 144788 3000
rect 144748 480 144776 2994
rect 145944 480 145972 4082
rect 146312 3738 146340 12022
rect 147692 3874 147720 12022
rect 147680 3868 147732 3874
rect 147680 3810 147732 3816
rect 146300 3732 146352 3738
rect 146300 3674 146352 3680
rect 148324 3732 148376 3738
rect 148324 3674 148376 3680
rect 147128 2984 147180 2990
rect 147128 2926 147180 2932
rect 147140 480 147168 2926
rect 148336 480 148364 3674
rect 149072 3466 149100 12022
rect 149060 3460 149112 3466
rect 149060 3402 149112 3408
rect 149520 3460 149572 3466
rect 149520 3402 149572 3408
rect 149532 480 149560 3402
rect 150452 3330 150480 12022
rect 150636 6914 150664 12022
rect 150544 6886 150664 6914
rect 150440 3324 150492 3330
rect 150440 3266 150492 3272
rect 150544 3058 150572 6886
rect 151832 4146 151860 12022
rect 151820 4140 151872 4146
rect 151820 4082 151872 4088
rect 150624 3868 150676 3874
rect 150624 3810 150676 3816
rect 150532 3052 150584 3058
rect 150532 2994 150584 3000
rect 150636 480 150664 3810
rect 151820 3528 151872 3534
rect 151820 3470 151872 3476
rect 151832 480 151860 3470
rect 153212 2990 153240 12022
rect 154592 3738 154620 12022
rect 156018 11778 156046 12036
rect 156800 12022 157136 12050
rect 157352 12022 158240 12050
rect 158732 12022 159344 12050
rect 160204 12022 160448 12050
rect 156018 11750 156092 11778
rect 155960 9512 156012 9518
rect 155960 9454 156012 9460
rect 155408 4072 155460 4078
rect 155408 4014 155460 4020
rect 154580 3732 154632 3738
rect 154580 3674 154632 3680
rect 154212 3324 154264 3330
rect 154212 3266 154264 3272
rect 153200 2984 153252 2990
rect 153200 2926 153252 2932
rect 153016 2916 153068 2922
rect 153016 2858 153068 2864
rect 153028 480 153056 2858
rect 154224 480 154252 3266
rect 155420 480 155448 4014
rect 155972 3874 156000 9454
rect 155960 3868 156012 3874
rect 155960 3810 156012 3816
rect 156064 3466 156092 11750
rect 156800 9518 156828 12022
rect 156788 9512 156840 9518
rect 156788 9454 156840 9460
rect 157352 3534 157380 12022
rect 157800 4140 157852 4146
rect 157800 4082 157852 4088
rect 157340 3528 157392 3534
rect 157340 3470 157392 3476
rect 156052 3460 156104 3466
rect 156052 3402 156104 3408
rect 156604 2984 156656 2990
rect 156604 2926 156656 2932
rect 156616 480 156644 2926
rect 157812 480 157840 4082
rect 158732 2922 158760 12022
rect 160100 3732 160152 3738
rect 160100 3674 160152 3680
rect 158904 3664 158956 3670
rect 158904 3606 158956 3612
rect 158720 2916 158772 2922
rect 158720 2858 158772 2864
rect 158916 480 158944 3606
rect 160112 480 160140 3674
rect 160204 3330 160232 12022
rect 161538 11778 161566 12036
rect 162320 12022 162656 12050
rect 162872 12022 163760 12050
rect 164252 12022 164864 12050
rect 165632 12022 165968 12050
rect 161538 11750 161612 11778
rect 161480 9512 161532 9518
rect 161480 9454 161532 9460
rect 161296 3460 161348 3466
rect 161296 3402 161348 3408
rect 160192 3324 160244 3330
rect 160192 3266 160244 3272
rect 161308 480 161336 3402
rect 161492 2990 161520 9454
rect 161584 4078 161612 11750
rect 162320 9518 162348 12022
rect 162308 9512 162360 9518
rect 162308 9454 162360 9460
rect 162872 4146 162900 12022
rect 162860 4140 162912 4146
rect 162860 4082 162912 4088
rect 161572 4072 161624 4078
rect 161572 4014 161624 4020
rect 163688 3800 163740 3806
rect 163688 3742 163740 3748
rect 162492 3324 162544 3330
rect 162492 3266 162544 3272
rect 161480 2984 161532 2990
rect 161480 2926 161532 2932
rect 162504 480 162532 3266
rect 163700 480 163728 3742
rect 164252 3670 164280 12022
rect 165632 3738 165660 12022
rect 167058 11778 167086 12036
rect 167840 12022 168176 12050
rect 168392 12022 169280 12050
rect 169772 12022 170384 12050
rect 171152 12022 171488 12050
rect 167058 11750 167132 11778
rect 167000 9512 167052 9518
rect 167000 9454 167052 9460
rect 166080 4004 166132 4010
rect 166080 3946 166132 3952
rect 165620 3732 165672 3738
rect 165620 3674 165672 3680
rect 164240 3664 164292 3670
rect 164240 3606 164292 3612
rect 164884 3256 164936 3262
rect 164884 3198 164936 3204
rect 164896 480 164924 3198
rect 166092 480 166120 3946
rect 167012 3330 167040 9454
rect 167104 3466 167132 11750
rect 167840 9518 167868 12022
rect 167828 9512 167880 9518
rect 167828 9454 167880 9460
rect 167184 3868 167236 3874
rect 167184 3810 167236 3816
rect 167092 3460 167144 3466
rect 167092 3402 167144 3408
rect 167000 3324 167052 3330
rect 167000 3266 167052 3272
rect 167196 480 167224 3810
rect 168392 3806 168420 12022
rect 168380 3800 168432 3806
rect 168380 3742 168432 3748
rect 169576 3664 169628 3670
rect 169576 3606 169628 3612
rect 168380 3528 168432 3534
rect 168380 3470 168432 3476
rect 168392 480 168420 3470
rect 169588 480 169616 3606
rect 169772 3262 169800 12022
rect 171152 4010 171180 12022
rect 172578 11778 172606 12036
rect 173360 12022 173696 12050
rect 173912 12022 174800 12050
rect 175292 12022 175904 12050
rect 176672 12022 177008 12050
rect 178052 12022 178112 12050
rect 178420 12022 179216 12050
rect 179432 12022 180320 12050
rect 180812 12022 181424 12050
rect 182192 12022 182528 12050
rect 183572 12022 183632 12050
rect 183940 12022 184736 12050
rect 184952 12022 185840 12050
rect 186332 12022 186944 12050
rect 187712 12022 188048 12050
rect 189092 12022 189152 12050
rect 189276 12022 190256 12050
rect 190472 12022 191360 12050
rect 191944 12022 192464 12050
rect 193324 12022 193568 12050
rect 194672 12022 194824 12050
rect 172578 11750 172652 11778
rect 172520 9512 172572 9518
rect 172520 9454 172572 9460
rect 171140 4004 171192 4010
rect 171140 3946 171192 3952
rect 171968 3732 172020 3738
rect 171968 3674 172020 3680
rect 170772 3596 170824 3602
rect 170772 3538 170824 3544
rect 169760 3256 169812 3262
rect 169760 3198 169812 3204
rect 170784 480 170812 3538
rect 171980 480 172008 3674
rect 172532 3534 172560 9454
rect 172624 3874 172652 11750
rect 173360 9518 173388 12022
rect 173348 9512 173400 9518
rect 173348 9454 173400 9460
rect 172612 3868 172664 3874
rect 172612 3810 172664 3816
rect 173912 3670 173940 12022
rect 173900 3664 173952 3670
rect 173900 3606 173952 3612
rect 175292 3602 175320 12022
rect 176672 3738 176700 12022
rect 177856 4072 177908 4078
rect 177856 4014 177908 4020
rect 176660 3732 176712 3738
rect 176660 3674 176712 3680
rect 175280 3596 175332 3602
rect 175280 3538 175332 3544
rect 172520 3528 172572 3534
rect 172520 3470 172572 3476
rect 174268 3528 174320 3534
rect 174268 3470 174320 3476
rect 173164 3188 173216 3194
rect 173164 3130 173216 3136
rect 173176 480 173204 3130
rect 174280 480 174308 3470
rect 175464 3460 175516 3466
rect 175464 3402 175516 3408
rect 175476 480 175504 3402
rect 176660 3324 176712 3330
rect 176660 3266 176712 3272
rect 176672 480 176700 3266
rect 177868 480 177896 4014
rect 178052 3194 178080 12022
rect 178420 6914 178448 12022
rect 178144 6886 178448 6914
rect 178144 3534 178172 6886
rect 178132 3528 178184 3534
rect 178132 3470 178184 3476
rect 179052 3528 179104 3534
rect 179052 3470 179104 3476
rect 178040 3188 178092 3194
rect 178040 3130 178092 3136
rect 179064 480 179092 3470
rect 179432 3466 179460 12022
rect 180248 3596 180300 3602
rect 180248 3538 180300 3544
rect 179420 3460 179472 3466
rect 179420 3402 179472 3408
rect 180260 480 180288 3538
rect 180812 3330 180840 12022
rect 182192 4078 182220 12022
rect 182180 4072 182232 4078
rect 182180 4014 182232 4020
rect 183572 3534 183600 12022
rect 183940 6914 183968 12022
rect 183664 6886 183968 6914
rect 183664 3602 183692 6886
rect 183652 3596 183704 3602
rect 183652 3538 183704 3544
rect 183560 3528 183612 3534
rect 183560 3470 183612 3476
rect 183744 3528 183796 3534
rect 183744 3470 183796 3476
rect 181444 3460 181496 3466
rect 181444 3402 181496 3408
rect 180800 3324 180852 3330
rect 180800 3266 180852 3272
rect 181456 480 181484 3402
rect 182548 3188 182600 3194
rect 182548 3130 182600 3136
rect 182560 480 182588 3130
rect 183756 480 183784 3470
rect 184952 3466 184980 12022
rect 184940 3460 184992 3466
rect 184940 3402 184992 3408
rect 186136 3324 186188 3330
rect 186136 3266 186188 3272
rect 184940 3256 184992 3262
rect 184940 3198 184992 3204
rect 184952 480 184980 3198
rect 186148 480 186176 3266
rect 186332 3194 186360 12022
rect 187332 4072 187384 4078
rect 187332 4014 187384 4020
rect 186320 3188 186372 3194
rect 186320 3130 186372 3136
rect 187344 480 187372 4014
rect 187712 3534 187740 12022
rect 188528 3868 188580 3874
rect 188528 3810 188580 3816
rect 187700 3528 187752 3534
rect 187700 3470 187752 3476
rect 188540 480 188568 3810
rect 189092 3262 189120 12022
rect 189276 6914 189304 12022
rect 189184 6886 189304 6914
rect 189184 3330 189212 6886
rect 190472 4078 190500 12022
rect 190460 4072 190512 4078
rect 190460 4014 190512 4020
rect 191944 3874 191972 12022
rect 192024 9512 192076 9518
rect 192024 9454 192076 9460
rect 191932 3868 191984 3874
rect 191932 3810 191984 3816
rect 189724 3528 189776 3534
rect 189724 3470 189776 3476
rect 189172 3324 189224 3330
rect 189172 3266 189224 3272
rect 189080 3256 189132 3262
rect 189080 3198 189132 3204
rect 189736 480 189764 3470
rect 190828 3460 190880 3466
rect 190828 3402 190880 3408
rect 190840 480 190868 3402
rect 192036 480 192064 9454
rect 193220 9444 193272 9450
rect 193220 9386 193272 9392
rect 193232 480 193260 9386
rect 193324 3534 193352 12022
rect 193312 3528 193364 3534
rect 193312 3470 193364 3476
rect 194796 3466 194824 12022
rect 195440 12022 195776 12050
rect 196544 12022 196880 12050
rect 197464 12022 197984 12050
rect 198844 12022 199088 12050
rect 195440 9518 195468 12022
rect 195428 9512 195480 9518
rect 195428 9454 195480 9460
rect 196544 9450 196572 12022
rect 196532 9444 196584 9450
rect 196532 9386 196584 9392
rect 196808 4072 196860 4078
rect 196808 4014 196860 4020
rect 194784 3460 194836 3466
rect 194784 3402 194836 3408
rect 194416 3324 194468 3330
rect 194416 3266 194468 3272
rect 194428 480 194456 3266
rect 195612 3256 195664 3262
rect 195612 3198 195664 3204
rect 195624 480 195652 3198
rect 196820 480 196848 4014
rect 197464 3330 197492 12022
rect 197912 8356 197964 8362
rect 197912 8298 197964 8304
rect 197452 3324 197504 3330
rect 197452 3266 197504 3272
rect 197924 480 197952 8298
rect 198844 3262 198872 12022
rect 200178 11778 200206 12036
rect 200960 12022 201296 12050
rect 202064 12022 202400 12050
rect 203168 12022 203504 12050
rect 204272 12022 204608 12050
rect 200178 11750 200252 11778
rect 199108 9240 199160 9246
rect 199108 9182 199160 9188
rect 198832 3256 198884 3262
rect 198832 3198 198884 3204
rect 199120 480 199148 9182
rect 200224 4078 200252 11750
rect 200304 9512 200356 9518
rect 200304 9454 200356 9460
rect 200212 4072 200264 4078
rect 200212 4014 200264 4020
rect 200316 480 200344 9454
rect 200960 8362 200988 12022
rect 202064 9246 202092 12022
rect 203168 9518 203196 12022
rect 203892 9580 203944 9586
rect 203892 9522 203944 9528
rect 203156 9512 203208 9518
rect 203156 9454 203208 9460
rect 202052 9240 202104 9246
rect 202052 9182 202104 9188
rect 201500 9172 201552 9178
rect 201500 9114 201552 9120
rect 200948 8356 201000 8362
rect 200948 8298 201000 8304
rect 201512 480 201540 9114
rect 202696 3324 202748 3330
rect 202696 3266 202748 3272
rect 202708 480 202736 3266
rect 203904 480 203932 9522
rect 204272 9178 204300 12022
rect 205698 11778 205726 12036
rect 206480 12022 206816 12050
rect 207584 12022 207920 12050
rect 208688 12022 209024 12050
rect 209884 12022 210128 12050
rect 211172 12022 211232 12050
rect 212000 12022 212336 12050
rect 213104 12022 213440 12050
rect 214208 12022 214544 12050
rect 215312 12022 215648 12050
rect 216692 12022 216752 12050
rect 217520 12022 217856 12050
rect 218624 12022 218960 12050
rect 219728 12022 220064 12050
rect 220832 12022 221168 12050
rect 222212 12022 222272 12050
rect 223040 12022 223376 12050
rect 224144 12022 224480 12050
rect 225248 12022 225584 12050
rect 226444 12022 226688 12050
rect 227732 12022 227792 12050
rect 228560 12022 228896 12050
rect 229664 12022 230000 12050
rect 230768 12022 231104 12050
rect 231872 12022 232208 12050
rect 233252 12022 233312 12050
rect 233436 12022 234416 12050
rect 234632 12022 235520 12050
rect 236288 12022 236624 12050
rect 237392 12022 237728 12050
rect 238772 12022 238832 12050
rect 239324 12022 239936 12050
rect 240152 12022 241040 12050
rect 241716 12022 242144 12050
rect 242912 12022 243248 12050
rect 244292 12022 244352 12050
rect 245212 12022 245456 12050
rect 245948 12022 246560 12050
rect 247604 12022 247664 12050
rect 248432 12022 248768 12050
rect 249872 12022 250024 12050
rect 250976 12022 251128 12050
rect 252080 12022 252416 12050
rect 253184 12022 253520 12050
rect 205698 11750 205772 11778
rect 205088 9444 205140 9450
rect 205088 9386 205140 9392
rect 204260 9172 204312 9178
rect 204260 9114 204312 9120
rect 205100 480 205128 9386
rect 205744 3330 205772 11750
rect 206480 9586 206508 12022
rect 206468 9580 206520 9586
rect 206468 9522 206520 9528
rect 206192 9512 206244 9518
rect 206192 9454 206244 9460
rect 205732 3324 205784 3330
rect 205732 3266 205784 3272
rect 206204 480 206232 9454
rect 207584 9450 207612 12022
rect 208688 9518 208716 12022
rect 208676 9512 208728 9518
rect 208676 9454 208728 9460
rect 209780 9512 209832 9518
rect 209780 9454 209832 9460
rect 207572 9444 207624 9450
rect 207572 9386 207624 9392
rect 207388 8492 207440 8498
rect 207388 8434 207440 8440
rect 207400 480 207428 8434
rect 208584 8424 208636 8430
rect 208584 8366 208636 8372
rect 208596 480 208624 8366
rect 209792 480 209820 9454
rect 209884 8498 209912 12022
rect 210976 9172 211028 9178
rect 210976 9114 211028 9120
rect 209872 8492 209924 8498
rect 209872 8434 209924 8440
rect 210988 480 211016 9114
rect 211172 8430 211200 12022
rect 212000 9518 212028 12022
rect 211988 9512 212040 9518
rect 211988 9454 212040 9460
rect 213104 9178 213132 12022
rect 213368 9444 213420 9450
rect 213368 9386 213420 9392
rect 213092 9172 213144 9178
rect 213092 9114 213144 9120
rect 212172 9036 212224 9042
rect 212172 8978 212224 8984
rect 211160 8424 211212 8430
rect 211160 8366 211212 8372
rect 212184 480 212212 8978
rect 213380 480 213408 9386
rect 214208 9042 214236 12022
rect 214472 9512 214524 9518
rect 214472 9454 214524 9460
rect 214196 9036 214248 9042
rect 214196 8978 214248 8984
rect 214484 480 214512 9454
rect 215312 9450 215340 12022
rect 216692 9518 216720 12022
rect 216680 9512 216732 9518
rect 216680 9454 216732 9460
rect 216864 9512 216916 9518
rect 216864 9454 216916 9460
rect 215300 9444 215352 9450
rect 215300 9386 215352 9392
rect 215668 9444 215720 9450
rect 215668 9386 215720 9392
rect 215680 480 215708 9386
rect 216876 480 216904 9454
rect 217520 9450 217548 12022
rect 218624 9518 218652 12022
rect 218612 9512 218664 9518
rect 218612 9454 218664 9460
rect 217508 9444 217560 9450
rect 217508 9386 217560 9392
rect 219256 8424 219308 8430
rect 219256 8366 219308 8372
rect 218060 8356 218112 8362
rect 218060 8298 218112 8304
rect 218072 480 218100 8298
rect 219268 480 219296 8366
rect 219728 8362 219756 12022
rect 220452 9512 220504 9518
rect 220452 9454 220504 9460
rect 219716 8356 219768 8362
rect 219716 8298 219768 8304
rect 220464 480 220492 9454
rect 220832 8430 220860 12022
rect 222212 9518 222240 12022
rect 222200 9512 222252 9518
rect 222200 9454 222252 9460
rect 222752 9512 222804 9518
rect 222752 9454 222804 9460
rect 221556 9444 221608 9450
rect 221556 9386 221608 9392
rect 220820 8424 220872 8430
rect 220820 8366 220872 8372
rect 221568 480 221596 9386
rect 222764 480 222792 9454
rect 223040 9450 223068 12022
rect 224144 9518 224172 12022
rect 224132 9512 224184 9518
rect 224132 9454 224184 9460
rect 223028 9444 223080 9450
rect 223028 9386 223080 9392
rect 225144 9444 225196 9450
rect 225144 9386 225196 9392
rect 223948 8764 224000 8770
rect 223948 8706 224000 8712
rect 223960 480 223988 8706
rect 225156 480 225184 9386
rect 225248 8770 225276 12022
rect 226340 9512 226392 9518
rect 226340 9454 226392 9460
rect 225236 8764 225288 8770
rect 225236 8706 225288 8712
rect 226352 480 226380 9454
rect 226444 9450 226472 12022
rect 227732 9518 227760 12022
rect 227720 9512 227772 9518
rect 227720 9454 227772 9460
rect 228560 9450 228588 12022
rect 228744 9654 229140 9674
rect 229664 9654 229692 12022
rect 228744 9648 229152 9654
rect 228744 9646 229100 9648
rect 226432 9444 226484 9450
rect 226432 9386 226484 9392
rect 227536 9444 227588 9450
rect 227536 9386 227588 9392
rect 228548 9444 228600 9450
rect 228548 9386 228600 9392
rect 227548 480 227576 9386
rect 228744 480 228772 9646
rect 229100 9590 229152 9596
rect 229652 9648 229704 9654
rect 229652 9590 229704 9596
rect 230768 8498 230796 12022
rect 231872 8770 231900 12022
rect 231032 8764 231084 8770
rect 231032 8706 231084 8712
rect 231860 8764 231912 8770
rect 231860 8706 231912 8712
rect 229836 8492 229888 8498
rect 229836 8434 229888 8440
rect 230756 8492 230808 8498
rect 230756 8434 230808 8440
rect 229848 480 229876 8434
rect 231044 480 231072 8706
rect 233252 8430 233280 12022
rect 232228 8424 232280 8430
rect 232228 8366 232280 8372
rect 233240 8424 233292 8430
rect 233240 8366 233292 8372
rect 232240 480 232268 8366
rect 233436 480 233464 12022
rect 234632 480 234660 12022
rect 236288 9518 236316 12022
rect 235816 9512 235868 9518
rect 235816 9454 235868 9460
rect 236276 9512 236328 9518
rect 237392 9466 237420 12022
rect 236276 9454 236328 9460
rect 235828 480 235856 9454
rect 237024 9438 237420 9466
rect 237024 480 237052 9438
rect 238772 8362 238800 12022
rect 238116 8356 238168 8362
rect 238116 8298 238168 8304
rect 238760 8356 238812 8362
rect 238760 8298 238812 8304
rect 238128 480 238156 8298
rect 239324 480 239352 12022
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240152 354 240180 12022
rect 241716 480 241744 12022
rect 242912 480 242940 12022
rect 244292 9466 244320 12022
rect 244108 9438 244320 9466
rect 244108 480 244136 9438
rect 245212 480 245240 12022
rect 240478 354 240590 480
rect 240152 326 240590 354
rect 240478 -960 240590 326
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 245948 354 245976 12022
rect 247604 480 247632 12022
rect 246366 354 246478 480
rect 245948 326 246478 354
rect 246366 -960 246478 326
rect 247562 -960 247674 480
rect 248432 354 248460 12022
rect 249996 480 250024 12022
rect 251100 9466 251128 12022
rect 251100 9438 251220 9466
rect 251192 480 251220 9438
rect 252388 480 252416 12022
rect 253492 480 253520 12022
rect 254228 12022 254288 12050
rect 255392 12022 255912 12050
rect 256496 12022 256648 12050
rect 257600 12022 257936 12050
rect 258704 12022 259040 12050
rect 248758 354 248870 480
rect 248432 326 248870 354
rect 248758 -960 248870 326
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254228 354 254256 12022
rect 255884 480 255912 12022
rect 256620 9518 256648 12022
rect 256608 9512 256660 9518
rect 256608 9454 256660 9460
rect 257068 9512 257120 9518
rect 257068 9454 257120 9460
rect 257080 480 257108 9454
rect 257908 8430 257936 12022
rect 259012 9518 259040 12022
rect 259472 12022 259808 12050
rect 260912 12022 261800 12050
rect 262016 12022 262168 12050
rect 263120 12022 263456 12050
rect 264224 12022 264560 12050
rect 265328 12022 265664 12050
rect 266432 12022 266768 12050
rect 267536 12022 267688 12050
rect 268640 12022 268976 12050
rect 269744 12022 270080 12050
rect 270848 12022 271184 12050
rect 271952 12022 272288 12050
rect 273056 12022 273208 12050
rect 274160 12022 274496 12050
rect 275264 12022 275600 12050
rect 276368 12022 276704 12050
rect 277472 12022 277808 12050
rect 278576 12022 278728 12050
rect 279680 12022 280016 12050
rect 280784 12022 281120 12050
rect 281888 12022 282224 12050
rect 282992 12022 283328 12050
rect 284096 12022 284248 12050
rect 285200 12022 285536 12050
rect 286304 12022 286640 12050
rect 287408 12022 287744 12050
rect 288512 12022 288848 12050
rect 289616 12022 289768 12050
rect 290720 12022 290964 12050
rect 291824 12022 292160 12050
rect 292928 12022 293264 12050
rect 294032 12022 294368 12050
rect 295136 12022 295288 12050
rect 296240 12022 296576 12050
rect 297344 12022 297680 12050
rect 298448 12022 298784 12050
rect 299552 12022 299888 12050
rect 300656 12022 300808 12050
rect 301760 12022 302096 12050
rect 302864 12022 303108 12050
rect 303968 12022 304304 12050
rect 305072 12022 305408 12050
rect 306176 12022 306328 12050
rect 307280 12022 307708 12050
rect 308384 12022 308720 12050
rect 309488 12022 309824 12050
rect 310592 12022 310928 12050
rect 311696 12022 311848 12050
rect 312800 12022 313136 12050
rect 313904 12022 314240 12050
rect 315008 12022 315344 12050
rect 316112 12022 316448 12050
rect 317216 12022 317368 12050
rect 318320 12022 318656 12050
rect 319424 12022 319760 12050
rect 320528 12022 320864 12050
rect 321632 12022 321968 12050
rect 322736 12022 322888 12050
rect 323840 12022 324084 12050
rect 324944 12022 325280 12050
rect 326048 12022 326384 12050
rect 327152 12022 327488 12050
rect 328256 12022 328408 12050
rect 329360 12022 329604 12050
rect 330464 12022 330800 12050
rect 331568 12022 331904 12050
rect 332672 12022 333008 12050
rect 333776 12022 333928 12050
rect 334880 12022 335216 12050
rect 335984 12022 336320 12050
rect 337088 12022 337424 12050
rect 338192 12022 338528 12050
rect 339296 12022 339448 12050
rect 340400 12022 340644 12050
rect 341504 12022 341840 12050
rect 342608 12022 342944 12050
rect 343712 12022 344048 12050
rect 344816 12022 344968 12050
rect 345920 12022 346348 12050
rect 347024 12022 347360 12050
rect 348128 12022 348464 12050
rect 349232 12022 349568 12050
rect 350336 12022 350488 12050
rect 351440 12022 351776 12050
rect 352544 12022 352880 12050
rect 353648 12022 353984 12050
rect 354752 12022 355088 12050
rect 355856 12022 356008 12050
rect 356960 12022 357296 12050
rect 358064 12022 358400 12050
rect 359168 12022 359504 12050
rect 360272 12022 360608 12050
rect 361376 12022 361528 12050
rect 362480 12022 362816 12050
rect 363584 12022 363920 12050
rect 364688 12022 365024 12050
rect 365792 12022 366128 12050
rect 366896 12022 367048 12050
rect 368000 12022 368244 12050
rect 369104 12022 369440 12050
rect 370208 12022 370544 12050
rect 371312 12022 371648 12050
rect 372416 12022 372568 12050
rect 373520 12022 373764 12050
rect 374624 12022 374960 12050
rect 375728 12022 376064 12050
rect 376832 12022 377168 12050
rect 259000 9512 259052 9518
rect 259000 9454 259052 9460
rect 257896 8424 257948 8430
rect 257896 8366 257948 8372
rect 258264 8424 258316 8430
rect 258264 8366 258316 8372
rect 258276 480 258304 8366
rect 259472 3602 259500 12022
rect 259552 9512 259604 9518
rect 259552 9454 259604 9460
rect 259460 3596 259512 3602
rect 259460 3538 259512 3544
rect 259564 3482 259592 9454
rect 260656 3596 260708 3602
rect 260656 3538 260708 3544
rect 259472 3454 259592 3482
rect 259472 480 259500 3454
rect 260668 480 260696 3538
rect 261772 480 261800 12022
rect 262140 9518 262168 12022
rect 262128 9512 262180 9518
rect 262128 9454 262180 9460
rect 262956 9512 263008 9518
rect 262956 9454 263008 9460
rect 262968 480 262996 9454
rect 263428 9178 263456 12022
rect 264532 9518 264560 12022
rect 264520 9512 264572 9518
rect 264520 9454 264572 9460
rect 265348 9512 265400 9518
rect 265348 9454 265400 9460
rect 263416 9172 263468 9178
rect 263416 9114 263468 9120
rect 264152 9172 264204 9178
rect 264152 9114 264204 9120
rect 264164 480 264192 9114
rect 265360 480 265388 9454
rect 265636 8906 265664 12022
rect 265624 8900 265676 8906
rect 265624 8842 265676 8848
rect 266544 8900 266596 8906
rect 266544 8842 266596 8848
rect 266556 480 266584 8842
rect 266740 8362 266768 12022
rect 267660 8566 267688 12022
rect 268948 9178 268976 12022
rect 270052 9518 270080 12022
rect 271156 9586 271184 12022
rect 271144 9580 271196 9586
rect 271144 9522 271196 9528
rect 270040 9512 270092 9518
rect 270040 9454 270092 9460
rect 271236 9512 271288 9518
rect 271236 9454 271288 9460
rect 268936 9172 268988 9178
rect 268936 9114 268988 9120
rect 270040 9172 270092 9178
rect 270040 9114 270092 9120
rect 267648 8560 267700 8566
rect 267648 8502 267700 8508
rect 268844 8560 268896 8566
rect 268844 8502 268896 8508
rect 266728 8356 266780 8362
rect 266728 8298 266780 8304
rect 267740 8356 267792 8362
rect 267740 8298 267792 8304
rect 267752 480 267780 8298
rect 268856 480 268884 8502
rect 270052 480 270080 9114
rect 271248 480 271276 9454
rect 272260 9450 272288 12022
rect 272432 9580 272484 9586
rect 272432 9522 272484 9528
rect 272248 9444 272300 9450
rect 272248 9386 272300 9392
rect 272444 480 272472 9522
rect 273180 9518 273208 12022
rect 273168 9512 273220 9518
rect 273168 9454 273220 9460
rect 274468 9450 274496 12022
rect 274548 9512 274600 9518
rect 274548 9454 274600 9460
rect 273628 9444 273680 9450
rect 273628 9386 273680 9392
rect 274456 9444 274508 9450
rect 274456 9386 274508 9392
rect 273640 480 273668 9386
rect 274560 3346 274588 9454
rect 275572 9246 275600 12022
rect 275928 9444 275980 9450
rect 275928 9386 275980 9392
rect 275560 9240 275612 9246
rect 275560 9182 275612 9188
rect 274560 3318 274864 3346
rect 274836 480 274864 3318
rect 275940 3074 275968 9386
rect 276676 8430 276704 12022
rect 277780 9518 277808 12022
rect 277768 9512 277820 9518
rect 277768 9454 277820 9460
rect 278700 9466 278728 12022
rect 279988 9518 280016 12022
rect 279516 9512 279568 9518
rect 278700 9438 278820 9466
rect 279516 9454 279568 9460
rect 279976 9512 280028 9518
rect 279976 9454 280028 9460
rect 277124 9240 277176 9246
rect 277124 9182 277176 9188
rect 276664 8424 276716 8430
rect 276664 8366 276716 8372
rect 275940 3046 276060 3074
rect 276032 480 276060 3046
rect 277136 480 277164 9182
rect 278320 8424 278372 8430
rect 278320 8366 278372 8372
rect 278332 480 278360 8366
rect 278792 3058 278820 9438
rect 278780 3052 278832 3058
rect 278780 2994 278832 3000
rect 279528 480 279556 9454
rect 281092 9450 281120 12022
rect 281448 9512 281500 9518
rect 281448 9454 281500 9460
rect 281080 9444 281132 9450
rect 281080 9386 281132 9392
rect 280712 3052 280764 3058
rect 280712 2994 280764 3000
rect 280724 480 280752 2994
rect 281460 2802 281488 9454
rect 282196 9382 282224 12022
rect 283300 9450 283328 12022
rect 284220 9518 284248 12022
rect 284208 9512 284260 9518
rect 284208 9454 284260 9460
rect 284668 9512 284720 9518
rect 284668 9454 284720 9460
rect 282828 9444 282880 9450
rect 282828 9386 282880 9392
rect 283288 9444 283340 9450
rect 283288 9386 283340 9392
rect 282184 9376 282236 9382
rect 282184 9318 282236 9324
rect 282840 3482 282868 9386
rect 284208 9376 284260 9382
rect 284208 9318 284260 9324
rect 284220 3482 284248 9318
rect 282840 3454 283144 3482
rect 284220 3454 284340 3482
rect 281460 2774 281580 2802
rect 254646 354 254758 480
rect 254228 326 254758 354
rect 254646 -960 254758 326
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281552 354 281580 2774
rect 283116 480 283144 3454
rect 284312 480 284340 3454
rect 284680 3058 284708 9454
rect 285404 9444 285456 9450
rect 285404 9386 285456 9392
rect 284668 3052 284720 3058
rect 284668 2994 284720 3000
rect 285416 480 285444 9386
rect 285508 8906 285536 12022
rect 285496 8900 285548 8906
rect 285496 8842 285548 8848
rect 286048 8900 286100 8906
rect 286048 8842 286100 8848
rect 286060 3874 286088 8842
rect 286612 8362 286640 12022
rect 287716 9518 287744 12022
rect 287704 9512 287756 9518
rect 287704 9454 287756 9460
rect 288440 9512 288492 9518
rect 288440 9454 288492 9460
rect 286600 8356 286652 8362
rect 286600 8298 286652 8304
rect 287244 8356 287296 8362
rect 287244 8298 287296 8304
rect 286048 3868 286100 3874
rect 286048 3810 286100 3816
rect 286600 3052 286652 3058
rect 286600 2994 286652 3000
rect 286612 480 286640 2994
rect 287256 2990 287284 8298
rect 287796 3868 287848 3874
rect 287796 3810 287848 3816
rect 287244 2984 287296 2990
rect 287244 2926 287296 2932
rect 287808 480 287836 3810
rect 288452 3058 288480 9454
rect 288820 8906 288848 12022
rect 289740 9450 289768 12022
rect 290936 9518 290964 12022
rect 290924 9512 290976 9518
rect 290924 9454 290976 9460
rect 291660 9512 291712 9518
rect 291660 9454 291712 9460
rect 289728 9444 289780 9450
rect 289728 9386 289780 9392
rect 291016 9444 291068 9450
rect 291016 9386 291068 9392
rect 288808 8900 288860 8906
rect 288808 8842 288860 8848
rect 291028 3534 291056 9386
rect 291108 8900 291160 8906
rect 291108 8842 291160 8848
rect 291016 3528 291068 3534
rect 291016 3470 291068 3476
rect 291120 3346 291148 8842
rect 291120 3318 291424 3346
rect 288440 3052 288492 3058
rect 288440 2994 288492 3000
rect 290188 3052 290240 3058
rect 290188 2994 290240 3000
rect 288992 2984 289044 2990
rect 288992 2926 289044 2932
rect 289004 480 289032 2926
rect 290200 480 290228 2994
rect 291396 480 291424 3318
rect 291672 3194 291700 9454
rect 292132 9450 292160 12022
rect 293236 9518 293264 12022
rect 293224 9512 293276 9518
rect 293224 9454 293276 9460
rect 294236 9512 294288 9518
rect 294236 9454 294288 9460
rect 292120 9444 292172 9450
rect 292120 9386 292172 9392
rect 292948 9444 293000 9450
rect 292948 9386 293000 9392
rect 292960 3534 292988 9386
rect 292580 3528 292632 3534
rect 292580 3470 292632 3476
rect 292948 3528 293000 3534
rect 292948 3470 293000 3476
rect 291660 3188 291712 3194
rect 291660 3130 291712 3136
rect 292592 480 292620 3470
rect 293684 3188 293736 3194
rect 293684 3130 293736 3136
rect 293696 480 293724 3130
rect 294248 3058 294276 9454
rect 294340 9450 294368 12022
rect 295260 9518 295288 12022
rect 295248 9512 295300 9518
rect 295248 9454 295300 9460
rect 296260 9512 296312 9518
rect 296260 9454 296312 9460
rect 294328 9444 294380 9450
rect 294328 9386 294380 9392
rect 295524 9444 295576 9450
rect 295524 9386 295576 9392
rect 295536 3874 295564 9386
rect 296272 4146 296300 9454
rect 296548 8362 296576 12022
rect 297652 9518 297680 12022
rect 297640 9512 297692 9518
rect 297640 9454 297692 9460
rect 298100 9512 298152 9518
rect 298100 9454 298152 9460
rect 296536 8356 296588 8362
rect 296536 8298 296588 8304
rect 296720 8356 296772 8362
rect 296720 8298 296772 8304
rect 296260 4140 296312 4146
rect 296260 4082 296312 4088
rect 295524 3868 295576 3874
rect 295524 3810 295576 3816
rect 294880 3528 294932 3534
rect 294880 3470 294932 3476
rect 294236 3052 294288 3058
rect 294236 2994 294288 3000
rect 294892 480 294920 3470
rect 296732 3330 296760 8298
rect 297272 3868 297324 3874
rect 297272 3810 297324 3816
rect 296720 3324 296772 3330
rect 296720 3266 296772 3272
rect 296076 3052 296128 3058
rect 296076 2994 296128 3000
rect 296088 480 296116 2994
rect 297284 480 297312 3810
rect 298112 3194 298140 9454
rect 298756 9178 298784 12022
rect 299860 9518 299888 12022
rect 299848 9512 299900 9518
rect 299848 9454 299900 9460
rect 300780 9450 300808 12022
rect 301320 9512 301372 9518
rect 301320 9454 301372 9460
rect 300768 9444 300820 9450
rect 300768 9386 300820 9392
rect 298744 9172 298796 9178
rect 298744 9114 298796 9120
rect 300676 9172 300728 9178
rect 300676 9114 300728 9120
rect 298468 4140 298520 4146
rect 298468 4082 298520 4088
rect 298100 3188 298152 3194
rect 298100 3130 298152 3136
rect 298480 480 298508 4082
rect 300688 3534 300716 9114
rect 300676 3528 300728 3534
rect 300676 3470 300728 3476
rect 301332 3466 301360 9454
rect 302068 9450 302096 12022
rect 303080 9518 303108 12022
rect 303068 9512 303120 9518
rect 303068 9454 303120 9460
rect 301872 9444 301924 9450
rect 301872 9386 301924 9392
rect 302056 9444 302108 9450
rect 302056 9386 302108 9392
rect 303160 9444 303212 9450
rect 303160 9386 303212 9392
rect 301320 3460 301372 3466
rect 301320 3402 301372 3408
rect 301884 3398 301912 9386
rect 303172 3602 303200 9386
rect 304276 9314 304304 12022
rect 304448 9512 304500 9518
rect 304448 9454 304500 9460
rect 304264 9308 304316 9314
rect 304264 9250 304316 9256
rect 304460 3738 304488 9454
rect 305380 8362 305408 12022
rect 305736 9308 305788 9314
rect 305736 9250 305788 9256
rect 305368 8356 305420 8362
rect 305368 8298 305420 8304
rect 305748 3874 305776 9250
rect 306300 8566 306328 12022
rect 307680 9466 307708 12022
rect 308692 9518 308720 12022
rect 308680 9512 308732 9518
rect 307680 9438 307800 9466
rect 308680 9454 308732 9460
rect 309796 9450 309824 12022
rect 310428 9512 310480 9518
rect 310428 9454 310480 9460
rect 306288 8560 306340 8566
rect 306288 8502 306340 8508
rect 306472 8560 306524 8566
rect 306472 8502 306524 8508
rect 305736 3868 305788 3874
rect 305736 3810 305788 3816
rect 304448 3732 304500 3738
rect 304448 3674 304500 3680
rect 303160 3596 303212 3602
rect 303160 3538 303212 3544
rect 305552 3596 305604 3602
rect 305552 3538 305604 3544
rect 301964 3528 302016 3534
rect 301964 3470 302016 3476
rect 301872 3392 301924 3398
rect 301872 3334 301924 3340
rect 299664 3324 299716 3330
rect 299664 3266 299716 3272
rect 299676 480 299704 3266
rect 300768 3188 300820 3194
rect 300768 3130 300820 3136
rect 300780 480 300808 3130
rect 301976 480 302004 3470
rect 303160 3460 303212 3466
rect 303160 3402 303212 3408
rect 303172 480 303200 3402
rect 304356 3392 304408 3398
rect 304356 3334 304408 3340
rect 304368 480 304396 3334
rect 305564 480 305592 3538
rect 306484 3330 306512 8502
rect 306932 8356 306984 8362
rect 306932 8298 306984 8304
rect 306748 3732 306800 3738
rect 306748 3674 306800 3680
rect 306472 3324 306524 3330
rect 306472 3266 306524 3272
rect 306760 480 306788 3674
rect 306944 3534 306972 8298
rect 306932 3528 306984 3534
rect 306932 3470 306984 3476
rect 307772 3466 307800 9438
rect 309784 9444 309836 9450
rect 309784 9386 309836 9392
rect 307944 3868 307996 3874
rect 307944 3810 307996 3816
rect 307760 3460 307812 3466
rect 307760 3402 307812 3408
rect 307956 480 307984 3810
rect 310440 3534 310468 9454
rect 310900 8498 310928 12022
rect 311820 9518 311848 12022
rect 311808 9512 311860 9518
rect 311808 9454 311860 9460
rect 311532 9444 311584 9450
rect 311532 9386 311584 9392
rect 310888 8492 310940 8498
rect 310888 8434 310940 8440
rect 309048 3528 309100 3534
rect 309048 3470 309100 3476
rect 310428 3528 310480 3534
rect 310428 3470 310480 3476
rect 309060 480 309088 3470
rect 311544 3466 311572 9386
rect 313108 8906 313136 12022
rect 314212 9518 314240 12022
rect 313188 9512 313240 9518
rect 313188 9454 313240 9460
rect 314200 9512 314252 9518
rect 314200 9454 314252 9460
rect 313096 8900 313148 8906
rect 313096 8842 313148 8848
rect 312728 8492 312780 8498
rect 312728 8434 312780 8440
rect 312636 3528 312688 3534
rect 312636 3470 312688 3476
rect 311440 3460 311492 3466
rect 311440 3402 311492 3408
rect 311532 3460 311584 3466
rect 311532 3402 311584 3408
rect 310244 3324 310296 3330
rect 310244 3266 310296 3272
rect 310256 480 310284 3266
rect 311452 480 311480 3402
rect 312648 480 312676 3470
rect 312740 3194 312768 8434
rect 313200 4010 313228 9454
rect 314568 8900 314620 8906
rect 314568 8842 314620 8848
rect 313188 4004 313240 4010
rect 313188 3946 313240 3952
rect 313832 3460 313884 3466
rect 313832 3402 313884 3408
rect 312728 3188 312780 3194
rect 312728 3130 312780 3136
rect 313844 480 313872 3402
rect 314580 3330 314608 8842
rect 315316 8566 315344 12022
rect 315856 9512 315908 9518
rect 315856 9454 315908 9460
rect 315304 8560 315356 8566
rect 315304 8502 315356 8508
rect 315868 3874 315896 9454
rect 316420 9382 316448 12022
rect 317340 9466 317368 12022
rect 317340 9438 317552 9466
rect 316408 9376 316460 9382
rect 316408 9318 316460 9324
rect 317420 9376 317472 9382
rect 317420 9318 317472 9324
rect 316040 8560 316092 8566
rect 316040 8502 316092 8508
rect 315856 3868 315908 3874
rect 315856 3810 315908 3816
rect 316052 3534 316080 8502
rect 316224 4004 316276 4010
rect 316224 3946 316276 3952
rect 316040 3528 316092 3534
rect 316040 3470 316092 3476
rect 314568 3324 314620 3330
rect 314568 3266 314620 3272
rect 315028 3188 315080 3194
rect 315028 3130 315080 3136
rect 315040 480 315068 3130
rect 316236 480 316264 3946
rect 317432 3330 317460 9318
rect 317524 3466 317552 9438
rect 318628 9178 318656 12022
rect 319732 9518 319760 12022
rect 319720 9512 319772 9518
rect 319720 9454 319772 9460
rect 320836 9382 320864 12022
rect 321940 9586 321968 12022
rect 321928 9580 321980 9586
rect 321928 9522 321980 9528
rect 322860 9518 322888 12022
rect 321468 9512 321520 9518
rect 321468 9454 321520 9460
rect 322848 9512 322900 9518
rect 322848 9454 322900 9460
rect 320824 9376 320876 9382
rect 320824 9318 320876 9324
rect 318616 9172 318668 9178
rect 318616 9114 318668 9120
rect 320088 9172 320140 9178
rect 320088 9114 320140 9120
rect 318524 3868 318576 3874
rect 318524 3810 318576 3816
rect 317512 3460 317564 3466
rect 317512 3402 317564 3408
rect 317328 3324 317380 3330
rect 317328 3266 317380 3272
rect 317420 3324 317472 3330
rect 317420 3266 317472 3272
rect 317340 480 317368 3266
rect 318536 480 318564 3810
rect 319720 3528 319772 3534
rect 319720 3470 319772 3476
rect 319732 480 319760 3470
rect 320100 3262 320128 9114
rect 320916 3324 320968 3330
rect 320916 3266 320968 3272
rect 320088 3256 320140 3262
rect 320088 3198 320140 3204
rect 320928 480 320956 3266
rect 321480 3194 321508 9454
rect 324056 9450 324084 12022
rect 324228 9580 324280 9586
rect 324228 9522 324280 9528
rect 324136 9512 324188 9518
rect 324136 9454 324188 9460
rect 324044 9444 324096 9450
rect 324044 9386 324096 9392
rect 322848 9376 322900 9382
rect 322848 9318 322900 9324
rect 322860 3534 322888 9318
rect 324148 4010 324176 9454
rect 324240 4146 324268 9522
rect 325252 9518 325280 12022
rect 325240 9512 325292 9518
rect 325240 9454 325292 9460
rect 326252 9512 326304 9518
rect 326252 9454 326304 9460
rect 325056 9444 325108 9450
rect 325056 9386 325108 9392
rect 324228 4140 324280 4146
rect 324228 4082 324280 4088
rect 324136 4004 324188 4010
rect 324136 3946 324188 3952
rect 322848 3528 322900 3534
rect 322848 3470 322900 3476
rect 325068 3466 325096 9386
rect 325608 3528 325660 3534
rect 325608 3470 325660 3476
rect 322112 3460 322164 3466
rect 322112 3402 322164 3408
rect 325056 3460 325108 3466
rect 325056 3402 325108 3408
rect 321468 3188 321520 3194
rect 321468 3130 321520 3136
rect 322124 480 322152 3402
rect 323308 3256 323360 3262
rect 323308 3198 323360 3204
rect 323320 480 323348 3198
rect 324412 3188 324464 3194
rect 324412 3130 324464 3136
rect 324424 480 324452 3130
rect 325620 480 325648 3470
rect 326264 3330 326292 9454
rect 326356 9450 326384 12022
rect 327460 9518 327488 12022
rect 327448 9512 327500 9518
rect 327448 9454 327500 9460
rect 328380 9450 328408 12022
rect 326344 9444 326396 9450
rect 326344 9386 326396 9392
rect 327080 9444 327132 9450
rect 327080 9386 327132 9392
rect 328368 9444 328420 9450
rect 328368 9386 328420 9392
rect 326804 4140 326856 4146
rect 326804 4082 326856 4088
rect 326252 3324 326304 3330
rect 326252 3266 326304 3272
rect 326816 480 326844 4082
rect 327092 3194 327120 9386
rect 329576 9178 329604 12022
rect 330772 9518 330800 12022
rect 329748 9512 329800 9518
rect 329748 9454 329800 9460
rect 330760 9512 330812 9518
rect 330760 9454 330812 9460
rect 329656 9444 329708 9450
rect 329656 9386 329708 9392
rect 329564 9172 329616 9178
rect 329564 9114 329616 9120
rect 328000 4004 328052 4010
rect 328000 3946 328052 3952
rect 327080 3188 327132 3194
rect 327080 3130 327132 3136
rect 328012 480 328040 3946
rect 329668 3466 329696 9386
rect 329760 3534 329788 9454
rect 331876 9382 331904 12022
rect 332508 9512 332560 9518
rect 332508 9454 332560 9460
rect 331864 9376 331916 9382
rect 331864 9318 331916 9324
rect 331128 9172 331180 9178
rect 331128 9114 331180 9120
rect 329748 3528 329800 3534
rect 329748 3470 329800 3476
rect 329196 3460 329248 3466
rect 329196 3402 329248 3408
rect 329656 3460 329708 3466
rect 329656 3402 329708 3408
rect 329208 480 329236 3402
rect 331140 3330 331168 9114
rect 332520 3942 332548 9454
rect 332980 9246 333008 12022
rect 333900 9466 333928 12022
rect 333900 9438 334296 9466
rect 333888 9376 333940 9382
rect 333888 9318 333940 9324
rect 332968 9240 333020 9246
rect 332968 9182 333020 9188
rect 333900 4146 333928 9318
rect 333888 4140 333940 4146
rect 333888 4082 333940 4088
rect 332508 3936 332560 3942
rect 332508 3878 332560 3884
rect 334268 3534 334296 9438
rect 335084 9240 335136 9246
rect 335084 9182 335136 9188
rect 335096 6914 335124 9182
rect 335188 8362 335216 12022
rect 336292 9518 336320 12022
rect 336280 9512 336332 9518
rect 336280 9454 336332 9460
rect 336740 9512 336792 9518
rect 336740 9454 336792 9460
rect 335176 8356 335228 8362
rect 335176 8298 335228 8304
rect 335360 8356 335412 8362
rect 335360 8298 335412 8304
rect 335096 6886 335216 6914
rect 335188 3806 335216 6886
rect 335176 3800 335228 3806
rect 335176 3742 335228 3748
rect 332692 3528 332744 3534
rect 332692 3470 332744 3476
rect 334256 3528 334308 3534
rect 334256 3470 334308 3476
rect 330392 3324 330444 3330
rect 330392 3266 330444 3272
rect 331128 3324 331180 3330
rect 331128 3266 331180 3272
rect 330404 480 330432 3266
rect 331588 3188 331640 3194
rect 331588 3130 331640 3136
rect 331600 480 331628 3130
rect 332704 480 332732 3470
rect 333888 3460 333940 3466
rect 333888 3402 333940 3408
rect 333900 480 333928 3402
rect 335372 3398 335400 8298
rect 336280 3936 336332 3942
rect 336280 3878 336332 3884
rect 335360 3392 335412 3398
rect 335360 3334 335412 3340
rect 335084 3324 335136 3330
rect 335084 3266 335136 3272
rect 335096 480 335124 3266
rect 336292 480 336320 3878
rect 336752 2922 336780 9454
rect 337396 9382 337424 12022
rect 338500 9586 338528 12022
rect 338488 9580 338540 9586
rect 338488 9522 338540 9528
rect 339420 9518 339448 12022
rect 339408 9512 339460 9518
rect 339408 9454 339460 9460
rect 340616 9450 340644 12022
rect 340788 9580 340840 9586
rect 340788 9522 340840 9528
rect 340696 9512 340748 9518
rect 340696 9454 340748 9460
rect 340604 9444 340656 9450
rect 340604 9386 340656 9392
rect 337384 9376 337436 9382
rect 337384 9318 337436 9324
rect 339408 9376 339460 9382
rect 339408 9318 339460 9324
rect 337476 4140 337528 4146
rect 337476 4082 337528 4088
rect 336740 2916 336792 2922
rect 336740 2858 336792 2864
rect 337488 480 337516 4082
rect 338672 3800 338724 3806
rect 338672 3742 338724 3748
rect 338684 480 338712 3742
rect 339420 3330 339448 9318
rect 340708 4078 340736 9454
rect 340696 4072 340748 4078
rect 340696 4014 340748 4020
rect 339868 3528 339920 3534
rect 339868 3470 339920 3476
rect 339408 3324 339460 3330
rect 339408 3266 339460 3272
rect 339880 480 339908 3470
rect 340800 3262 340828 9522
rect 341812 9518 341840 12022
rect 341800 9512 341852 9518
rect 341800 9454 341852 9460
rect 342168 9444 342220 9450
rect 342168 9386 342220 9392
rect 342180 4146 342208 9386
rect 342916 9314 342944 12022
rect 343548 9512 343600 9518
rect 343548 9454 343600 9460
rect 342904 9308 342956 9314
rect 342904 9250 342956 9256
rect 342168 4140 342220 4146
rect 342168 4082 342220 4088
rect 343560 3534 343588 9454
rect 343732 9308 343784 9314
rect 343732 9250 343784 9256
rect 343548 3528 343600 3534
rect 343548 3470 343600 3476
rect 343744 3466 343772 9250
rect 344020 8702 344048 12022
rect 344940 9246 344968 12022
rect 346320 9466 346348 12022
rect 347332 9518 347360 12022
rect 347320 9512 347372 9518
rect 346320 9438 346440 9466
rect 347320 9454 347372 9460
rect 344928 9240 344980 9246
rect 344928 9182 344980 9188
rect 345112 9240 345164 9246
rect 345112 9182 345164 9188
rect 344008 8696 344060 8702
rect 344008 8638 344060 8644
rect 345020 8696 345072 8702
rect 345020 8638 345072 8644
rect 343732 3460 343784 3466
rect 343732 3402 343784 3408
rect 340972 3392 341024 3398
rect 340972 3334 341024 3340
rect 340788 3256 340840 3262
rect 340788 3198 340840 3204
rect 340984 480 341012 3334
rect 345032 3330 345060 8638
rect 345124 3398 345152 9182
rect 345756 4072 345808 4078
rect 345756 4014 345808 4020
rect 345112 3392 345164 3398
rect 345112 3334 345164 3340
rect 343364 3324 343416 3330
rect 343364 3266 343416 3272
rect 345020 3324 345072 3330
rect 345020 3266 345072 3272
rect 342168 2916 342220 2922
rect 342168 2858 342220 2864
rect 342180 480 342208 2858
rect 343376 480 343404 3266
rect 344560 3256 344612 3262
rect 344560 3198 344612 3204
rect 344572 480 344600 3198
rect 345768 480 345796 4014
rect 346412 3602 346440 9438
rect 348436 8634 348464 12022
rect 349068 9512 349120 9518
rect 349068 9454 349120 9460
rect 348424 8628 348476 8634
rect 348424 8570 348476 8576
rect 346952 4140 347004 4146
rect 346952 4082 347004 4088
rect 346400 3596 346452 3602
rect 346400 3538 346452 3544
rect 346964 480 346992 4082
rect 348056 3528 348108 3534
rect 348056 3470 348108 3476
rect 348068 480 348096 3470
rect 349080 2922 349108 9454
rect 349540 9450 349568 12022
rect 350460 9518 350488 12022
rect 351748 9518 351776 12022
rect 350448 9512 350500 9518
rect 350448 9454 350500 9460
rect 351092 9512 351144 9518
rect 351092 9454 351144 9460
rect 351736 9512 351788 9518
rect 351736 9454 351788 9460
rect 349528 9444 349580 9450
rect 349528 9386 349580 9392
rect 350448 8628 350500 8634
rect 350448 8570 350500 8576
rect 350460 4078 350488 8570
rect 350448 4072 350500 4078
rect 350448 4014 350500 4020
rect 351104 3466 351132 9454
rect 352852 9450 352880 12022
rect 353208 9512 353260 9518
rect 353208 9454 353260 9460
rect 351828 9444 351880 9450
rect 351828 9386 351880 9392
rect 352840 9444 352892 9450
rect 352840 9386 352892 9392
rect 351840 4146 351868 9386
rect 351828 4140 351880 4146
rect 351828 4082 351880 4088
rect 353220 3670 353248 9454
rect 353956 8974 353984 12022
rect 355060 9518 355088 12022
rect 355048 9512 355100 9518
rect 355048 9454 355100 9460
rect 355980 9466 356008 12022
rect 357268 9518 357296 12022
rect 356152 9512 356204 9518
rect 354496 9444 354548 9450
rect 355980 9438 356100 9466
rect 356152 9454 356204 9460
rect 357256 9512 357308 9518
rect 357256 9454 357308 9460
rect 354496 9386 354548 9392
rect 353944 8968 353996 8974
rect 353944 8910 353996 8916
rect 354508 3738 354536 9386
rect 355048 8968 355100 8974
rect 355048 8910 355100 8916
rect 354496 3732 354548 3738
rect 354496 3674 354548 3680
rect 353208 3664 353260 3670
rect 353208 3606 353260 3612
rect 352840 3596 352892 3602
rect 352840 3538 352892 3544
rect 349252 3460 349304 3466
rect 349252 3402 349304 3408
rect 351092 3460 351144 3466
rect 351092 3402 351144 3408
rect 349068 2916 349120 2922
rect 349068 2858 349120 2864
rect 349264 480 349292 3402
rect 351644 3392 351696 3398
rect 351644 3334 351696 3340
rect 350448 3324 350500 3330
rect 350448 3266 350500 3272
rect 350460 480 350488 3266
rect 351656 480 351684 3334
rect 352852 480 352880 3538
rect 355060 3534 355088 8910
rect 355232 4072 355284 4078
rect 355232 4014 355284 4020
rect 355048 3528 355100 3534
rect 355048 3470 355100 3476
rect 354036 2916 354088 2922
rect 354036 2858 354088 2864
rect 354048 480 354076 2858
rect 355244 480 355272 4014
rect 356072 3262 356100 9438
rect 356060 3256 356112 3262
rect 356060 3198 356112 3204
rect 356164 3058 356192 9454
rect 358372 9450 358400 12022
rect 358728 9512 358780 9518
rect 358728 9454 358780 9460
rect 358360 9444 358412 9450
rect 358360 9386 358412 9392
rect 358740 4146 358768 9454
rect 359476 9314 359504 12022
rect 360108 9444 360160 9450
rect 360108 9386 360160 9392
rect 359464 9308 359516 9314
rect 359464 9250 359516 9256
rect 356336 4140 356388 4146
rect 356336 4082 356388 4088
rect 358728 4140 358780 4146
rect 358728 4082 358780 4088
rect 356152 3052 356204 3058
rect 356152 2994 356204 3000
rect 356348 480 356376 4082
rect 360120 4010 360148 9386
rect 360580 8906 360608 12022
rect 361500 9450 361528 12022
rect 361488 9444 361540 9450
rect 361488 9386 361540 9392
rect 361488 9308 361540 9314
rect 361488 9250 361540 9256
rect 360568 8900 360620 8906
rect 360568 8842 360620 8848
rect 361500 4078 361528 9250
rect 362788 9042 362816 12022
rect 362868 9444 362920 9450
rect 362868 9386 362920 9392
rect 362776 9036 362828 9042
rect 362776 8978 362828 8984
rect 362776 8900 362828 8906
rect 362776 8842 362828 8848
rect 361488 4072 361540 4078
rect 361488 4014 361540 4020
rect 360108 4004 360160 4010
rect 360108 3946 360160 3952
rect 362788 3874 362816 8842
rect 362776 3868 362828 3874
rect 362776 3810 362828 3816
rect 362880 3806 362908 9386
rect 363328 9036 363380 9042
rect 363328 8978 363380 8984
rect 362868 3800 362920 3806
rect 362868 3742 362920 3748
rect 359924 3732 359976 3738
rect 359924 3674 359976 3680
rect 358728 3664 358780 3670
rect 358728 3606 358780 3612
rect 357532 3460 357584 3466
rect 357532 3402 357584 3408
rect 357544 480 357572 3402
rect 358740 480 358768 3606
rect 359936 480 359964 3674
rect 363340 3670 363368 8978
rect 363892 8838 363920 12022
rect 364996 9042 365024 12022
rect 366100 9518 366128 12022
rect 366088 9512 366140 9518
rect 366088 9454 366140 9460
rect 367020 9450 367048 12022
rect 367008 9444 367060 9450
rect 367008 9386 367060 9392
rect 364984 9036 365036 9042
rect 364984 8978 365036 8984
rect 365720 9036 365772 9042
rect 365720 8978 365772 8984
rect 363880 8832 363932 8838
rect 363880 8774 363932 8780
rect 364800 8832 364852 8838
rect 364800 8774 364852 8780
rect 364616 4140 364668 4146
rect 364616 4082 364668 4088
rect 363328 3664 363380 3670
rect 363328 3606 363380 3612
rect 361120 3528 361172 3534
rect 361120 3470 361172 3476
rect 361132 480 361160 3470
rect 363512 3256 363564 3262
rect 363512 3198 363564 3204
rect 362316 3052 362368 3058
rect 362316 2994 362368 3000
rect 362328 480 362356 2994
rect 363524 480 363552 3198
rect 364628 480 364656 4082
rect 364812 3058 364840 8774
rect 365732 3466 365760 8978
rect 368216 8634 368244 12022
rect 368388 9512 368440 9518
rect 368388 9454 368440 9460
rect 368296 9444 368348 9450
rect 368296 9386 368348 9392
rect 368204 8628 368256 8634
rect 368204 8570 368256 8576
rect 368308 4146 368336 9386
rect 368296 4140 368348 4146
rect 368296 4082 368348 4088
rect 367008 4072 367060 4078
rect 367008 4014 367060 4020
rect 365812 4004 365864 4010
rect 365812 3946 365864 3952
rect 365720 3460 365772 3466
rect 365720 3402 365772 3408
rect 364800 3052 364852 3058
rect 364800 2994 364852 3000
rect 365824 480 365852 3946
rect 367020 480 367048 4014
rect 368204 3868 368256 3874
rect 368204 3810 368256 3816
rect 368216 480 368244 3810
rect 368400 3602 368428 9454
rect 369412 9450 369440 12022
rect 370516 9518 370544 12022
rect 370504 9512 370556 9518
rect 370504 9454 370556 9460
rect 369400 9444 369452 9450
rect 369400 9386 369452 9392
rect 371148 9444 371200 9450
rect 371148 9386 371200 9392
rect 369768 8628 369820 8634
rect 369768 8570 369820 8576
rect 369780 4078 369808 8570
rect 369768 4072 369820 4078
rect 369768 4014 369820 4020
rect 369400 3800 369452 3806
rect 369400 3742 369452 3748
rect 368388 3596 368440 3602
rect 368388 3538 368440 3544
rect 369412 480 369440 3742
rect 371160 3670 371188 9386
rect 371620 9042 371648 12022
rect 372540 9518 372568 12022
rect 372160 9512 372212 9518
rect 372160 9454 372212 9460
rect 372528 9512 372580 9518
rect 372528 9454 372580 9460
rect 373356 9512 373408 9518
rect 373356 9454 373408 9460
rect 371608 9036 371660 9042
rect 371608 8978 371660 8984
rect 372172 3806 372200 9454
rect 372620 9036 372672 9042
rect 372620 8978 372672 8984
rect 372632 3942 372660 8978
rect 372620 3936 372672 3942
rect 372620 3878 372672 3884
rect 372160 3800 372212 3806
rect 372160 3742 372212 3748
rect 370596 3664 370648 3670
rect 370596 3606 370648 3612
rect 371148 3664 371200 3670
rect 371148 3606 371200 3612
rect 370608 480 370636 3606
rect 373368 3466 373396 9454
rect 373736 9110 373764 12022
rect 374932 9450 374960 12022
rect 376036 9518 376064 12022
rect 376024 9512 376076 9518
rect 376024 9454 376076 9460
rect 374920 9444 374972 9450
rect 374920 9386 374972 9392
rect 375380 9444 375432 9450
rect 375380 9386 375432 9392
rect 373724 9104 373776 9110
rect 373724 9046 373776 9052
rect 374368 9104 374420 9110
rect 374368 9046 374420 9052
rect 374092 3596 374144 3602
rect 374092 3538 374144 3544
rect 372896 3460 372948 3466
rect 372896 3402 372948 3408
rect 373356 3460 373408 3466
rect 373356 3402 373408 3408
rect 371700 3052 371752 3058
rect 371700 2994 371752 3000
rect 371712 480 371740 2994
rect 372908 480 372936 3402
rect 374104 480 374132 3538
rect 374380 3126 374408 9046
rect 375288 4140 375340 4146
rect 375288 4082 375340 4088
rect 374368 3120 374420 3126
rect 374368 3062 374420 3068
rect 375300 480 375328 4082
rect 375392 2990 375420 9386
rect 377140 9110 377168 12022
rect 377876 12022 377936 12050
rect 379040 12022 379376 12050
rect 380144 12022 380480 12050
rect 381248 12022 381584 12050
rect 382352 12022 382688 12050
rect 383456 12022 383608 12050
rect 384560 12022 384988 12050
rect 385664 12022 386000 12050
rect 386768 12022 387104 12050
rect 387872 12022 388208 12050
rect 388976 12022 389128 12050
rect 390080 12022 390416 12050
rect 391184 12022 391520 12050
rect 392288 12022 392624 12050
rect 393392 12022 393728 12050
rect 394496 12022 394648 12050
rect 395600 12022 396028 12050
rect 396704 12022 397040 12050
rect 397808 12022 398144 12050
rect 398912 12022 399248 12050
rect 400016 12022 400168 12050
rect 401120 12022 401364 12050
rect 402224 12022 402560 12050
rect 403328 12022 403664 12050
rect 404432 12022 404768 12050
rect 405536 12022 405688 12050
rect 406640 12022 406976 12050
rect 407744 12022 408080 12050
rect 408848 12022 409184 12050
rect 409952 12022 410288 12050
rect 377876 9382 377904 12022
rect 378048 9512 378100 9518
rect 378048 9454 378100 9460
rect 377864 9376 377916 9382
rect 377864 9318 377916 9324
rect 377128 9104 377180 9110
rect 377128 9046 377180 9052
rect 376484 4072 376536 4078
rect 376484 4014 376536 4020
rect 375380 2984 375432 2990
rect 375380 2926 375432 2932
rect 376496 480 376524 4014
rect 378060 4010 378088 9454
rect 379244 9104 379296 9110
rect 379244 9046 379296 9052
rect 379256 6914 379284 9046
rect 379348 8430 379376 12022
rect 380452 9518 380480 12022
rect 381556 9586 381584 12022
rect 381544 9580 381596 9586
rect 381544 9522 381596 9528
rect 380440 9512 380492 9518
rect 380440 9454 380492 9460
rect 381728 9512 381780 9518
rect 381728 9454 381780 9460
rect 379428 9376 379480 9382
rect 379428 9318 379480 9324
rect 379336 8424 379388 8430
rect 379336 8366 379388 8372
rect 379256 6886 379376 6914
rect 378048 4004 378100 4010
rect 378048 3946 378100 3952
rect 378876 3800 378928 3806
rect 378876 3742 378928 3748
rect 377680 3664 377732 3670
rect 377680 3606 377732 3612
rect 377692 480 377720 3606
rect 378888 480 378916 3742
rect 379348 3330 379376 6886
rect 379440 3806 379468 9318
rect 380808 8424 380860 8430
rect 380808 8366 380860 8372
rect 379980 3936 380032 3942
rect 379980 3878 380032 3884
rect 379428 3800 379480 3806
rect 379428 3742 379480 3748
rect 379336 3324 379388 3330
rect 379336 3266 379388 3272
rect 379992 480 380020 3878
rect 380820 3602 380848 8366
rect 380808 3596 380860 3602
rect 380808 3538 380860 3544
rect 381740 3466 381768 9454
rect 382660 9246 382688 12022
rect 382924 9580 382976 9586
rect 382924 9522 382976 9528
rect 382648 9240 382700 9246
rect 382648 9182 382700 9188
rect 382936 3738 382964 9522
rect 383580 8566 383608 12022
rect 384960 9466 384988 12022
rect 385972 9518 386000 12022
rect 385960 9512 386012 9518
rect 384960 9438 385080 9466
rect 385960 9454 386012 9460
rect 384396 9240 384448 9246
rect 384396 9182 384448 9188
rect 383568 8560 383620 8566
rect 383568 8502 383620 8508
rect 383660 8560 383712 8566
rect 383660 8502 383712 8508
rect 382924 3732 382976 3738
rect 382924 3674 382976 3680
rect 381176 3460 381228 3466
rect 381176 3402 381228 3408
rect 381728 3460 381780 3466
rect 381728 3402 381780 3408
rect 381188 480 381216 3402
rect 382372 3120 382424 3126
rect 382372 3062 382424 3068
rect 382384 480 382412 3062
rect 383672 3058 383700 8502
rect 383660 3052 383712 3058
rect 383660 2994 383712 3000
rect 384408 2990 384436 9182
rect 384764 4004 384816 4010
rect 384764 3946 384816 3952
rect 383568 2984 383620 2990
rect 383568 2926 383620 2932
rect 384396 2984 384448 2990
rect 384396 2926 384448 2932
rect 383580 480 383608 2926
rect 384776 480 384804 3946
rect 385052 3670 385080 9438
rect 387076 9382 387104 12022
rect 387708 9512 387760 9518
rect 387708 9454 387760 9460
rect 387064 9376 387116 9382
rect 387064 9318 387116 9324
rect 387720 4146 387748 9454
rect 388180 8906 388208 12022
rect 389100 9518 389128 12022
rect 389088 9512 389140 9518
rect 389088 9454 389140 9460
rect 390388 9450 390416 12022
rect 391492 9518 391520 12022
rect 390468 9512 390520 9518
rect 390468 9454 390520 9460
rect 391480 9512 391532 9518
rect 391480 9454 391532 9460
rect 392492 9512 392544 9518
rect 392492 9454 392544 9460
rect 390376 9444 390428 9450
rect 390376 9386 390428 9392
rect 389088 9376 389140 9382
rect 389088 9318 389140 9324
rect 388168 8900 388220 8906
rect 388168 8842 388220 8848
rect 387708 4140 387760 4146
rect 387708 4082 387760 4088
rect 389100 4010 389128 9318
rect 390192 8900 390244 8906
rect 390192 8842 390244 8848
rect 389088 4004 389140 4010
rect 389088 3946 389140 3952
rect 387156 3800 387208 3806
rect 387156 3742 387208 3748
rect 385040 3664 385092 3670
rect 385040 3606 385092 3612
rect 385960 3324 386012 3330
rect 385960 3266 386012 3272
rect 385972 480 386000 3266
rect 387168 480 387196 3742
rect 388260 3596 388312 3602
rect 388260 3538 388312 3544
rect 388272 480 388300 3538
rect 390204 3466 390232 8842
rect 390480 3534 390508 9454
rect 391848 9444 391900 9450
rect 391848 9386 391900 9392
rect 391860 3806 391888 9386
rect 392504 3942 392532 9454
rect 392596 8566 392624 12022
rect 393700 9382 393728 12022
rect 394620 9466 394648 12022
rect 396000 9466 396028 12022
rect 397012 9518 397040 12022
rect 397000 9512 397052 9518
rect 394620 9438 394924 9466
rect 396000 9438 396304 9466
rect 397000 9454 397052 9460
rect 393688 9376 393740 9382
rect 393688 9318 393740 9324
rect 394792 9376 394844 9382
rect 394792 9318 394844 9324
rect 392584 8560 392636 8566
rect 392584 8502 392636 8508
rect 393320 8560 393372 8566
rect 393320 8502 393372 8508
rect 392492 3936 392544 3942
rect 392492 3878 392544 3884
rect 391848 3800 391900 3806
rect 391848 3742 391900 3748
rect 390652 3732 390704 3738
rect 390652 3674 390704 3680
rect 390468 3528 390520 3534
rect 390468 3470 390520 3476
rect 389456 3460 389508 3466
rect 389456 3402 389508 3408
rect 390192 3460 390244 3466
rect 390192 3402 390244 3408
rect 389468 480 389496 3402
rect 390664 480 390692 3674
rect 393332 3398 393360 8502
rect 394804 3874 394832 9318
rect 394792 3868 394844 3874
rect 394792 3810 394844 3816
rect 394896 3738 394924 9438
rect 395344 4140 395396 4146
rect 395344 4082 395396 4088
rect 394884 3732 394936 3738
rect 394884 3674 394936 3680
rect 394240 3596 394292 3602
rect 394240 3538 394292 3544
rect 393320 3392 393372 3398
rect 393320 3334 393372 3340
rect 393044 3052 393096 3058
rect 393044 2994 393096 3000
rect 391848 2984 391900 2990
rect 391848 2926 391900 2932
rect 391860 480 391888 2926
rect 393056 480 393084 2994
rect 394252 480 394280 3538
rect 395356 480 395384 4082
rect 396276 3602 396304 9438
rect 398116 9382 398144 12022
rect 398748 9512 398800 9518
rect 398748 9454 398800 9460
rect 398104 9376 398156 9382
rect 398104 9318 398156 9324
rect 396540 4004 396592 4010
rect 396540 3946 396592 3952
rect 396264 3596 396316 3602
rect 396264 3538 396316 3544
rect 396552 480 396580 3946
rect 398760 3466 398788 9454
rect 399220 8906 399248 12022
rect 400140 9518 400168 12022
rect 400128 9512 400180 9518
rect 400128 9454 400180 9460
rect 401336 9450 401364 12022
rect 401416 9512 401468 9518
rect 401416 9454 401468 9460
rect 401324 9444 401376 9450
rect 401324 9386 401376 9392
rect 400128 9376 400180 9382
rect 400128 9318 400180 9324
rect 399208 8900 399260 8906
rect 399208 8842 399260 8848
rect 400140 3806 400168 9318
rect 401428 3942 401456 9454
rect 402532 8974 402560 12022
rect 402888 9444 402940 9450
rect 402888 9386 402940 9392
rect 402520 8968 402572 8974
rect 402520 8910 402572 8916
rect 401508 8900 401560 8906
rect 401508 8842 401560 8848
rect 401520 4010 401548 8842
rect 401508 4004 401560 4010
rect 401508 3946 401560 3952
rect 401324 3936 401376 3942
rect 401324 3878 401376 3884
rect 401416 3936 401468 3942
rect 401416 3878 401468 3884
rect 400036 3800 400088 3806
rect 400036 3742 400088 3748
rect 400128 3800 400180 3806
rect 400128 3742 400180 3748
rect 398932 3528 398984 3534
rect 398932 3470 398984 3476
rect 397736 3460 397788 3466
rect 397736 3402 397788 3408
rect 398748 3460 398800 3466
rect 398748 3402 398800 3408
rect 397748 480 397776 3402
rect 398944 480 398972 3470
rect 400048 1986 400076 3742
rect 400048 1958 400168 1986
rect 400140 480 400168 1958
rect 401336 480 401364 3878
rect 402900 3670 402928 9386
rect 403636 9314 403664 12022
rect 403624 9308 403676 9314
rect 403624 9250 403676 9256
rect 404360 9308 404412 9314
rect 404360 9250 404412 9256
rect 403440 8968 403492 8974
rect 403440 8910 403492 8916
rect 402888 3664 402940 3670
rect 402888 3606 402940 3612
rect 403452 3602 403480 8910
rect 403624 3868 403676 3874
rect 403624 3810 403676 3816
rect 403440 3596 403492 3602
rect 403440 3538 403492 3544
rect 402520 3392 402572 3398
rect 402520 3334 402572 3340
rect 402532 480 402560 3334
rect 403636 480 403664 3810
rect 404372 3398 404400 9250
rect 404740 8770 404768 12022
rect 405660 9450 405688 12022
rect 406948 9518 406976 12022
rect 408052 9518 408080 12022
rect 409156 9518 409184 12022
rect 410260 9586 410288 12022
rect 410996 12022 411056 12050
rect 412160 12022 412496 12050
rect 413264 12022 413600 12050
rect 414368 12022 414704 12050
rect 415472 12022 415808 12050
rect 410248 9580 410300 9586
rect 410248 9522 410300 9528
rect 406936 9512 406988 9518
rect 406936 9454 406988 9460
rect 407396 9512 407448 9518
rect 407396 9454 407448 9460
rect 408040 9512 408092 9518
rect 408040 9454 408092 9460
rect 408500 9512 408552 9518
rect 408500 9454 408552 9460
rect 409144 9512 409196 9518
rect 409144 9454 409196 9460
rect 405648 9444 405700 9450
rect 405648 9386 405700 9392
rect 407028 9444 407080 9450
rect 407028 9386 407080 9392
rect 404728 8764 404780 8770
rect 404728 8706 404780 8712
rect 406108 8764 406160 8770
rect 406108 8706 406160 8712
rect 406120 4078 406148 8706
rect 406108 4072 406160 4078
rect 406108 4014 406160 4020
rect 407040 3738 407068 9386
rect 407408 3874 407436 9454
rect 407396 3868 407448 3874
rect 407396 3810 407448 3816
rect 408408 3800 408460 3806
rect 408408 3742 408460 3748
rect 404820 3732 404872 3738
rect 404820 3674 404872 3680
rect 407028 3732 407080 3738
rect 407028 3674 407080 3680
rect 404360 3392 404412 3398
rect 404360 3334 404412 3340
rect 404832 480 404860 3674
rect 406016 3528 406068 3534
rect 406016 3470 406068 3476
rect 406028 480 406056 3470
rect 407212 3460 407264 3466
rect 407212 3402 407264 3408
rect 407224 480 407252 3402
rect 408420 480 408448 3742
rect 408512 3330 408540 9454
rect 410996 9450 411024 12022
rect 412364 9580 412416 9586
rect 412364 9522 412416 9528
rect 411168 9512 411220 9518
rect 411168 9454 411220 9460
rect 410984 9444 411036 9450
rect 410984 9386 411036 9392
rect 409604 4004 409656 4010
rect 409604 3946 409656 3952
rect 408500 3324 408552 3330
rect 408500 3266 408552 3272
rect 409616 480 409644 3946
rect 411180 3942 411208 9454
rect 412376 4010 412404 9522
rect 412468 8430 412496 12022
rect 413572 9518 413600 12022
rect 413560 9512 413612 9518
rect 413560 9454 413612 9460
rect 414020 9512 414072 9518
rect 414020 9454 414072 9460
rect 412548 9444 412600 9450
rect 412548 9386 412600 9392
rect 412456 8424 412508 8430
rect 412456 8366 412508 8372
rect 412364 4004 412416 4010
rect 412364 3946 412416 3952
rect 410800 3936 410852 3942
rect 410800 3878 410852 3884
rect 411168 3936 411220 3942
rect 411168 3878 411220 3884
rect 410812 480 410840 3878
rect 412560 3670 412588 9386
rect 412640 8424 412692 8430
rect 412640 8366 412692 8372
rect 411904 3664 411956 3670
rect 411904 3606 411956 3612
rect 412548 3664 412600 3670
rect 412548 3606 412600 3612
rect 411916 480 411944 3606
rect 412652 3534 412680 8366
rect 413100 3596 413152 3602
rect 413100 3538 413152 3544
rect 412640 3528 412692 3534
rect 412640 3470 412692 3476
rect 413112 480 413140 3538
rect 414032 3466 414060 9454
rect 414676 9450 414704 12022
rect 414664 9444 414716 9450
rect 414664 9386 414716 9392
rect 415780 9314 415808 12022
rect 416516 12022 416576 12050
rect 417680 12022 418016 12050
rect 418784 12022 419120 12050
rect 419888 12022 420224 12050
rect 420992 12022 421328 12050
rect 422096 12022 422248 12050
rect 423200 12022 423628 12050
rect 424304 12022 424640 12050
rect 425408 12022 425744 12050
rect 426512 12022 426848 12050
rect 416516 9518 416544 12022
rect 416504 9512 416556 9518
rect 416504 9454 416556 9460
rect 417988 9450 418016 12022
rect 419092 9518 419120 12022
rect 418068 9512 418120 9518
rect 418068 9454 418120 9460
rect 419080 9512 419132 9518
rect 419080 9454 419132 9460
rect 416688 9444 416740 9450
rect 416688 9386 416740 9392
rect 417976 9444 418028 9450
rect 417976 9386 418028 9392
rect 415768 9308 415820 9314
rect 415768 9250 415820 9256
rect 416700 4146 416728 9386
rect 417976 9308 418028 9314
rect 417976 9250 418028 9256
rect 416688 4140 416740 4146
rect 416688 4082 416740 4088
rect 415492 4072 415544 4078
rect 415492 4014 415544 4020
rect 414020 3460 414072 3466
rect 414020 3402 414072 3408
rect 414296 3392 414348 3398
rect 414296 3334 414348 3340
rect 414308 480 414336 3334
rect 415504 480 415532 4014
rect 417884 3868 417936 3874
rect 417884 3810 417936 3816
rect 416688 3732 416740 3738
rect 416688 3674 416740 3680
rect 416700 480 416728 3674
rect 417896 480 417924 3810
rect 417988 3398 418016 9250
rect 418080 3874 418108 9454
rect 419448 9444 419500 9450
rect 419448 9386 419500 9392
rect 418068 3868 418120 3874
rect 418068 3810 418120 3816
rect 419460 3466 419488 9386
rect 420196 8770 420224 12022
rect 420828 9512 420880 9518
rect 420828 9454 420880 9460
rect 420184 8764 420236 8770
rect 420184 8706 420236 8712
rect 420184 3936 420236 3942
rect 420184 3878 420236 3884
rect 419448 3460 419500 3466
rect 419448 3402 419500 3408
rect 417976 3392 418028 3398
rect 417976 3334 418028 3340
rect 418988 3324 419040 3330
rect 418988 3266 419040 3272
rect 419000 480 419028 3266
rect 420196 480 420224 3878
rect 420840 3806 420868 9454
rect 420920 8764 420972 8770
rect 420920 8706 420972 8712
rect 420828 3800 420880 3806
rect 420828 3742 420880 3748
rect 420932 3602 420960 8706
rect 421300 8566 421328 12022
rect 421288 8560 421340 8566
rect 421288 8502 421340 8508
rect 422220 8362 422248 12022
rect 423600 9466 423628 12022
rect 423600 9438 423812 9466
rect 423036 8560 423088 8566
rect 423036 8502 423088 8508
rect 422208 8356 422260 8362
rect 422208 8298 422260 8304
rect 422300 8356 422352 8362
rect 422300 8298 422352 8304
rect 422312 4010 422340 8298
rect 423048 4078 423076 8502
rect 423036 4072 423088 4078
rect 423036 4014 423088 4020
rect 421380 4004 421432 4010
rect 421380 3946 421432 3952
rect 422300 4004 422352 4010
rect 422300 3946 422352 3952
rect 420920 3596 420972 3602
rect 420920 3538 420972 3544
rect 421392 480 421420 3946
rect 423784 3738 423812 9438
rect 424612 8634 424640 12022
rect 425716 9178 425744 12022
rect 426820 9518 426848 12022
rect 427556 12022 427616 12050
rect 428720 12022 429056 12050
rect 429824 12022 430160 12050
rect 430928 12022 431264 12050
rect 432032 12022 432368 12050
rect 433136 12022 433288 12050
rect 434240 12022 434576 12050
rect 435344 12022 435680 12050
rect 436448 12022 436784 12050
rect 437552 12022 437888 12050
rect 438656 12022 438808 12050
rect 439760 12022 440096 12050
rect 440864 12022 441200 12050
rect 441968 12022 442304 12050
rect 443072 12022 443408 12050
rect 444176 12022 444328 12050
rect 445280 12022 445616 12050
rect 446384 12022 446720 12050
rect 447488 12022 447824 12050
rect 448592 12022 448928 12050
rect 449696 12022 449848 12050
rect 450800 12022 451136 12050
rect 451904 12022 452240 12050
rect 453008 12022 453252 12050
rect 454112 12022 454448 12050
rect 455216 12022 455368 12050
rect 456320 12022 456564 12050
rect 457424 12022 457760 12050
rect 458528 12022 458864 12050
rect 459632 12022 459968 12050
rect 460736 12022 460888 12050
rect 461840 12022 462176 12050
rect 462944 12022 463280 12050
rect 464048 12022 464384 12050
rect 465152 12022 465488 12050
rect 466256 12022 466408 12050
rect 467360 12022 467696 12050
rect 468464 12022 468800 12050
rect 469568 12022 469904 12050
rect 470672 12022 471008 12050
rect 426808 9512 426860 9518
rect 426808 9454 426860 9460
rect 425704 9172 425756 9178
rect 425704 9114 425756 9120
rect 427556 9110 427584 12022
rect 427820 9512 427872 9518
rect 427820 9454 427872 9460
rect 427728 9172 427780 9178
rect 427728 9114 427780 9120
rect 427544 9104 427596 9110
rect 427544 9046 427596 9052
rect 424600 8628 424652 8634
rect 424600 8570 424652 8576
rect 426072 8628 426124 8634
rect 426072 8570 426124 8576
rect 423772 3732 423824 3738
rect 423772 3674 423824 3680
rect 422576 3664 422628 3670
rect 422576 3606 422628 3612
rect 422588 480 422616 3606
rect 426084 3534 426112 8570
rect 426164 4140 426216 4146
rect 426164 4082 426216 4088
rect 423772 3528 423824 3534
rect 423772 3470 423824 3476
rect 426072 3528 426124 3534
rect 426072 3470 426124 3476
rect 423784 480 423812 3470
rect 424968 3392 425020 3398
rect 424968 3334 425020 3340
rect 424980 480 425008 3334
rect 426176 480 426204 4082
rect 427740 3942 427768 9114
rect 427728 3936 427780 3942
rect 427728 3878 427780 3884
rect 427832 3670 427860 9454
rect 429028 9314 429056 12022
rect 429016 9308 429068 9314
rect 429016 9250 429068 9256
rect 429660 9308 429712 9314
rect 429660 9250 429712 9256
rect 429672 3874 429700 9250
rect 430132 8566 430160 12022
rect 431236 8974 431264 12022
rect 432340 9450 432368 12022
rect 432328 9444 432380 9450
rect 432328 9386 432380 9392
rect 433260 9382 433288 12022
rect 433340 9444 433392 9450
rect 433340 9386 433392 9392
rect 433248 9376 433300 9382
rect 433248 9318 433300 9324
rect 431224 8968 431276 8974
rect 431224 8910 431276 8916
rect 432236 8968 432288 8974
rect 432236 8910 432288 8916
rect 430120 8560 430172 8566
rect 430120 8502 430172 8508
rect 430948 8560 431000 8566
rect 430948 8502 431000 8508
rect 428464 3868 428516 3874
rect 428464 3810 428516 3816
rect 429660 3868 429712 3874
rect 429660 3810 429712 3816
rect 427820 3664 427872 3670
rect 427820 3606 427872 3612
rect 427268 3324 427320 3330
rect 427268 3266 427320 3272
rect 427280 480 427308 3266
rect 428476 480 428504 3810
rect 430960 3806 430988 8502
rect 430856 3800 430908 3806
rect 430856 3742 430908 3748
rect 430948 3800 431000 3806
rect 430948 3742 431000 3748
rect 429660 3460 429712 3466
rect 429660 3402 429712 3408
rect 429672 480 429700 3402
rect 430868 480 430896 3742
rect 432248 3602 432276 8910
rect 433248 4072 433300 4078
rect 433248 4014 433300 4020
rect 432052 3596 432104 3602
rect 432052 3538 432104 3544
rect 432236 3596 432288 3602
rect 432236 3538 432288 3544
rect 432064 480 432092 3538
rect 433260 480 433288 4014
rect 433352 3466 433380 9386
rect 434548 8974 434576 12022
rect 435652 9042 435680 12022
rect 436756 9314 436784 12022
rect 437860 9450 437888 12022
rect 437848 9444 437900 9450
rect 437848 9386 437900 9392
rect 438780 9314 438808 12022
rect 438860 9444 438912 9450
rect 438860 9386 438912 9392
rect 436744 9308 436796 9314
rect 436744 9250 436796 9256
rect 438676 9308 438728 9314
rect 438676 9250 438728 9256
rect 438768 9308 438820 9314
rect 438768 9250 438820 9256
rect 435640 9036 435692 9042
rect 435640 8978 435692 8984
rect 434536 8968 434588 8974
rect 434536 8910 434588 8916
rect 434444 4004 434496 4010
rect 434444 3946 434496 3952
rect 433340 3460 433392 3466
rect 433340 3402 433392 3408
rect 434456 480 434484 3946
rect 437940 3936 437992 3942
rect 437940 3878 437992 3884
rect 435548 3732 435600 3738
rect 435548 3674 435600 3680
rect 435560 480 435588 3674
rect 436744 3528 436796 3534
rect 436744 3470 436796 3476
rect 436756 480 436784 3470
rect 437952 480 437980 3878
rect 438688 3738 438716 9250
rect 438676 3732 438728 3738
rect 438676 3674 438728 3680
rect 438872 3534 438900 9386
rect 440068 9178 440096 12022
rect 440056 9172 440108 9178
rect 440056 9114 440108 9120
rect 440332 9104 440384 9110
rect 440332 9046 440384 9052
rect 439136 3664 439188 3670
rect 439136 3606 439188 3612
rect 438860 3528 438912 3534
rect 438860 3470 438912 3476
rect 439148 480 439176 3606
rect 440344 480 440372 9046
rect 441172 8634 441200 12022
rect 442276 9246 442304 12022
rect 443380 9450 443408 12022
rect 444300 9518 444328 12022
rect 445588 9586 445616 12022
rect 445576 9580 445628 9586
rect 445576 9522 445628 9528
rect 444288 9512 444340 9518
rect 444288 9454 444340 9460
rect 443368 9444 443420 9450
rect 443368 9386 443420 9392
rect 446220 9376 446272 9382
rect 446220 9318 446272 9324
rect 442264 9240 442316 9246
rect 442264 9182 442316 9188
rect 441160 8628 441212 8634
rect 441160 8570 441212 8576
rect 441528 3868 441580 3874
rect 441528 3810 441580 3816
rect 441540 480 441568 3810
rect 442632 3800 442684 3806
rect 442632 3742 442684 3748
rect 442644 480 442672 3742
rect 443828 3596 443880 3602
rect 443828 3538 443880 3544
rect 443840 480 443868 3538
rect 445024 3460 445076 3466
rect 445024 3402 445076 3408
rect 445036 480 445064 3402
rect 446232 480 446260 9318
rect 446692 8838 446720 12022
rect 447796 9110 447824 12022
rect 448900 9654 448928 12022
rect 448888 9648 448940 9654
rect 448888 9590 448940 9596
rect 449820 9110 449848 12022
rect 447784 9104 447836 9110
rect 447784 9046 447836 9052
rect 449808 9104 449860 9110
rect 449808 9046 449860 9052
rect 448612 9036 448664 9042
rect 448612 8978 448664 8984
rect 447416 8968 447468 8974
rect 447416 8910 447468 8916
rect 446680 8832 446732 8838
rect 446680 8774 446732 8780
rect 447428 480 447456 8910
rect 448624 480 448652 8978
rect 451108 8974 451136 12022
rect 452108 9308 452160 9314
rect 452108 9250 452160 9256
rect 451096 8968 451148 8974
rect 451096 8910 451148 8916
rect 449808 3732 449860 3738
rect 449808 3674 449860 3680
rect 449820 480 449848 3674
rect 450912 3528 450964 3534
rect 450912 3470 450964 3476
rect 450924 480 450952 3470
rect 452120 480 452148 9250
rect 452212 8702 452240 12022
rect 453224 8770 453252 12022
rect 453304 9172 453356 9178
rect 453304 9114 453356 9120
rect 453212 8764 453264 8770
rect 453212 8706 453264 8712
rect 452200 8696 452252 8702
rect 452200 8638 452252 8644
rect 453316 480 453344 9114
rect 454420 8566 454448 12022
rect 455340 9314 455368 12022
rect 456536 9382 456564 12022
rect 457732 9450 457760 12022
rect 458088 9512 458140 9518
rect 458088 9454 458140 9460
rect 456892 9444 456944 9450
rect 456892 9386 456944 9392
rect 457720 9444 457772 9450
rect 457720 9386 457772 9392
rect 456524 9376 456576 9382
rect 456524 9318 456576 9324
rect 455328 9308 455380 9314
rect 455328 9250 455380 9256
rect 455696 9240 455748 9246
rect 455696 9182 455748 9188
rect 454500 8628 454552 8634
rect 454500 8570 454552 8576
rect 454408 8560 454460 8566
rect 454408 8502 454460 8508
rect 454512 480 454540 8570
rect 455708 480 455736 9182
rect 456904 480 456932 9386
rect 458100 480 458128 9454
rect 458836 9246 458864 12022
rect 459192 9580 459244 9586
rect 459192 9522 459244 9528
rect 458824 9240 458876 9246
rect 458824 9182 458876 9188
rect 459204 480 459232 9522
rect 459940 8498 459968 12022
rect 460860 8838 460888 12022
rect 462148 9042 462176 12022
rect 463252 9654 463280 12022
rect 462780 9648 462832 9654
rect 462780 9590 462832 9596
rect 463240 9648 463292 9654
rect 463240 9590 463292 9596
rect 462320 9172 462372 9178
rect 462320 9114 462372 9120
rect 461584 9036 461636 9042
rect 461584 8978 461636 8984
rect 462136 9036 462188 9042
rect 462136 8978 462188 8984
rect 460388 8832 460440 8838
rect 460388 8774 460440 8780
rect 460848 8832 460900 8838
rect 460848 8774 460900 8780
rect 459928 8492 459980 8498
rect 459928 8434 459980 8440
rect 460400 480 460428 8774
rect 461596 480 461624 8978
rect 462332 3534 462360 9114
rect 462320 3528 462372 3534
rect 462320 3470 462372 3476
rect 462792 480 462820 9590
rect 464356 9110 464384 12022
rect 465460 9178 465488 12022
rect 465448 9172 465500 9178
rect 465448 9114 465500 9120
rect 464344 9104 464396 9110
rect 464344 9046 464396 9052
rect 464988 8968 465040 8974
rect 464988 8910 465040 8916
rect 463976 3528 464028 3534
rect 463976 3470 464028 3476
rect 465000 3482 465028 8910
rect 466276 8696 466328 8702
rect 466276 8638 466328 8644
rect 463988 480 464016 3470
rect 465000 3454 465212 3482
rect 465184 480 465212 3454
rect 466288 480 466316 8638
rect 466380 8634 466408 12022
rect 467668 9586 467696 12022
rect 467656 9580 467708 9586
rect 467656 9522 467708 9528
rect 467840 9308 467892 9314
rect 467840 9250 467892 9256
rect 467472 8764 467524 8770
rect 467472 8706 467524 8712
rect 466368 8628 466420 8634
rect 466368 8570 466420 8576
rect 467484 480 467512 8706
rect 467852 3534 467880 9250
rect 468772 8702 468800 12022
rect 469876 9518 469904 12022
rect 469864 9512 469916 9518
rect 469864 9454 469916 9460
rect 470508 9376 470560 9382
rect 470508 9318 470560 9324
rect 468760 8696 468812 8702
rect 468760 8638 468812 8644
rect 468668 8560 468720 8566
rect 468668 8502 468720 8508
rect 467840 3528 467892 3534
rect 467840 3470 467892 3476
rect 468680 480 468708 8502
rect 469864 3528 469916 3534
rect 469864 3470 469916 3476
rect 469876 480 469904 3470
rect 470520 2802 470548 9318
rect 470980 8974 471008 12022
rect 471716 12022 471776 12050
rect 472880 12022 473216 12050
rect 473984 12022 474320 12050
rect 475088 12022 475424 12050
rect 476192 12022 476528 12050
rect 477296 12022 477448 12050
rect 478400 12022 478736 12050
rect 479504 12022 479840 12050
rect 480608 12022 480944 12050
rect 481712 12022 482048 12050
rect 482816 12022 482968 12050
rect 483920 12022 484256 12050
rect 485024 12022 485360 12050
rect 486128 12022 486464 12050
rect 487232 12022 487568 12050
rect 488336 12022 488488 12050
rect 489440 12022 489684 12050
rect 490544 12022 490880 12050
rect 491648 12022 491984 12050
rect 492752 12022 493088 12050
rect 470968 8968 471020 8974
rect 470968 8910 471020 8916
rect 471716 8906 471744 12022
rect 473188 9450 473216 12022
rect 471888 9444 471940 9450
rect 471888 9386 471940 9392
rect 473176 9444 473228 9450
rect 473176 9386 473228 9392
rect 471704 8900 471756 8906
rect 471704 8842 471756 8848
rect 471900 3482 471928 9386
rect 471980 9240 472032 9246
rect 471980 9182 472032 9188
rect 471992 3602 472020 9182
rect 474292 8770 474320 12022
rect 475396 9246 475424 12022
rect 476304 9648 476356 9654
rect 476304 9590 476356 9596
rect 475384 9240 475436 9246
rect 475384 9182 475436 9188
rect 475108 9036 475160 9042
rect 475108 8978 475160 8984
rect 474648 8832 474700 8838
rect 474648 8774 474700 8780
rect 474280 8764 474332 8770
rect 474280 8706 474332 8712
rect 474556 8492 474608 8498
rect 474556 8434 474608 8440
rect 471980 3596 472032 3602
rect 471980 3538 472032 3544
rect 473452 3596 473504 3602
rect 473452 3538 473504 3544
rect 471900 3454 472296 3482
rect 470520 2774 470640 2802
rect 281878 354 281990 480
rect 281552 326 281990 354
rect 281878 -960 281990 326
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 470612 354 470640 2774
rect 472268 480 472296 3454
rect 473464 480 473492 3538
rect 474568 480 474596 8434
rect 474660 3534 474688 8774
rect 474648 3528 474700 3534
rect 474648 3470 474700 3476
rect 475120 3058 475148 8978
rect 476316 3534 476344 9590
rect 476500 9382 476528 12022
rect 476488 9376 476540 9382
rect 476488 9318 476540 9324
rect 477420 9042 477448 12022
rect 478708 9654 478736 12022
rect 478696 9648 478748 9654
rect 478696 9590 478748 9596
rect 478788 9104 478840 9110
rect 478788 9046 478840 9052
rect 477408 9036 477460 9042
rect 477408 8978 477460 8984
rect 475752 3528 475804 3534
rect 475752 3470 475804 3476
rect 476304 3528 476356 3534
rect 476304 3470 476356 3476
rect 478144 3528 478196 3534
rect 478144 3470 478196 3476
rect 475108 3052 475160 3058
rect 475108 2994 475160 3000
rect 475764 480 475792 3470
rect 476948 3052 477000 3058
rect 476948 2994 477000 3000
rect 476960 480 476988 2994
rect 478156 480 478184 3470
rect 478800 2802 478828 9046
rect 479812 8838 479840 12022
rect 480628 9580 480680 9586
rect 480628 9522 480680 9528
rect 480168 9172 480220 9178
rect 480168 9114 480220 9120
rect 479800 8832 479852 8838
rect 479800 8774 479852 8780
rect 478880 8628 478932 8634
rect 478880 8570 478932 8576
rect 478892 3806 478920 8570
rect 480180 4026 480208 9114
rect 480180 3998 480576 4026
rect 478880 3800 478932 3806
rect 478880 3742 478932 3748
rect 478800 2774 478920 2802
rect 471030 354 471142 480
rect 470612 326 471142 354
rect 471030 -960 471142 326
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 478892 354 478920 2774
rect 480548 480 480576 3998
rect 480640 3534 480668 9522
rect 480916 9178 480944 12022
rect 482020 9314 482048 12022
rect 482940 9586 482968 12022
rect 482928 9580 482980 9586
rect 482928 9522 482980 9528
rect 482008 9308 482060 9314
rect 482008 9250 482060 9256
rect 480904 9172 480956 9178
rect 480904 9114 480956 9120
rect 484228 9110 484256 12022
rect 484308 9512 484360 9518
rect 484308 9454 484360 9460
rect 484216 9104 484268 9110
rect 484216 9046 484268 9052
rect 481640 8696 481692 8702
rect 481640 8638 481692 8644
rect 480628 3528 480680 3534
rect 480628 3470 480680 3476
rect 481652 3466 481680 8638
rect 481732 3800 481784 3806
rect 481732 3742 481784 3748
rect 481640 3460 481692 3466
rect 481640 3402 481692 3408
rect 481744 480 481772 3742
rect 484320 3534 484348 9454
rect 484676 8968 484728 8974
rect 484676 8910 484728 8916
rect 482836 3528 482888 3534
rect 482836 3470 482888 3476
rect 484308 3528 484360 3534
rect 484308 3470 484360 3476
rect 482848 480 482876 3470
rect 484032 3460 484084 3466
rect 484032 3402 484084 3408
rect 484044 480 484072 3402
rect 484688 2990 484716 8910
rect 485332 8702 485360 12022
rect 486436 9518 486464 12022
rect 486424 9512 486476 9518
rect 486424 9454 486476 9460
rect 486332 9444 486384 9450
rect 486332 9386 486384 9392
rect 485688 8900 485740 8906
rect 485688 8842 485740 8848
rect 485320 8696 485372 8702
rect 485320 8638 485372 8644
rect 485228 3528 485280 3534
rect 485228 3470 485280 3476
rect 484676 2984 484728 2990
rect 484676 2926 484728 2932
rect 485240 480 485268 3470
rect 485700 3058 485728 8842
rect 486344 3194 486372 9386
rect 487540 8974 487568 12022
rect 487528 8968 487580 8974
rect 487528 8910 487580 8916
rect 488460 8906 488488 12022
rect 489656 9450 489684 12022
rect 489644 9444 489696 9450
rect 489644 9386 489696 9392
rect 490104 9376 490156 9382
rect 490104 9318 490156 9324
rect 488540 9240 488592 9246
rect 488540 9182 488592 9188
rect 488448 8900 488500 8906
rect 488448 8842 488500 8848
rect 487160 8764 487212 8770
rect 487160 8706 487212 8712
rect 487172 3466 487200 8706
rect 488552 4010 488580 9182
rect 490012 9036 490064 9042
rect 490012 8978 490064 8984
rect 488540 4004 488592 4010
rect 488540 3946 488592 3952
rect 487160 3460 487212 3466
rect 487160 3402 487212 3408
rect 489920 3460 489972 3466
rect 489920 3402 489972 3408
rect 486332 3188 486384 3194
rect 486332 3130 486384 3136
rect 488816 3188 488868 3194
rect 488816 3130 488868 3136
rect 485688 3052 485740 3058
rect 485688 2994 485740 3000
rect 487620 3052 487672 3058
rect 487620 2994 487672 3000
rect 486424 2984 486476 2990
rect 486424 2926 486476 2932
rect 486436 480 486464 2926
rect 487632 480 487660 2994
rect 488828 480 488856 3130
rect 489932 480 489960 3402
rect 490024 3194 490052 8978
rect 490116 3534 490144 9318
rect 490852 9246 490880 12022
rect 491392 9648 491444 9654
rect 491392 9590 491444 9596
rect 490840 9240 490892 9246
rect 490840 9182 490892 9188
rect 491116 4004 491168 4010
rect 491116 3946 491168 3952
rect 490104 3528 490156 3534
rect 490104 3470 490156 3476
rect 490012 3188 490064 3194
rect 490012 3130 490064 3136
rect 491128 480 491156 3946
rect 491404 3602 491432 9590
rect 491956 8634 491984 12022
rect 493060 9042 493088 12022
rect 493796 12022 493856 12050
rect 494960 12022 495296 12050
rect 496064 12022 496400 12050
rect 497168 12022 497504 12050
rect 498272 12022 498608 12050
rect 499376 12022 499528 12050
rect 500480 12022 500816 12050
rect 501584 12022 501920 12050
rect 502688 12022 503024 12050
rect 503792 12022 504128 12050
rect 504896 12022 505048 12050
rect 506000 12022 506336 12050
rect 507104 12022 507440 12050
rect 508208 12022 508544 12050
rect 509312 12022 509648 12050
rect 510416 12022 510568 12050
rect 511520 12022 511856 12050
rect 512624 12022 512960 12050
rect 513728 12022 514064 12050
rect 514832 12022 515168 12050
rect 515936 12022 516088 12050
rect 517040 12022 517376 12050
rect 518144 12022 518480 12050
rect 519248 12022 519584 12050
rect 520352 12022 520688 12050
rect 521456 12022 521608 12050
rect 522560 12022 522896 12050
rect 523664 12022 524000 12050
rect 524768 12022 525104 12050
rect 493048 9036 493100 9042
rect 493048 8978 493100 8984
rect 491944 8628 491996 8634
rect 491944 8570 491996 8576
rect 493796 8498 493824 12022
rect 493968 8832 494020 8838
rect 493968 8774 494020 8780
rect 493784 8492 493836 8498
rect 493784 8434 493836 8440
rect 491392 3596 491444 3602
rect 491392 3538 491444 3544
rect 492312 3528 492364 3534
rect 492312 3470 492364 3476
rect 492324 480 492352 3470
rect 493508 3188 493560 3194
rect 493508 3130 493560 3136
rect 493520 480 493548 3130
rect 493980 3058 494008 8774
rect 495268 8770 495296 12022
rect 496372 9382 496400 12022
rect 496452 9580 496504 9586
rect 496452 9522 496504 9528
rect 496360 9376 496412 9382
rect 496360 9318 496412 9324
rect 495532 9308 495584 9314
rect 495532 9250 495584 9256
rect 495348 9172 495400 9178
rect 495348 9114 495400 9120
rect 495256 8764 495308 8770
rect 495256 8706 495308 8712
rect 494704 3596 494756 3602
rect 494704 3538 494756 3544
rect 493968 3052 494020 3058
rect 493968 2994 494020 3000
rect 494716 480 494744 3538
rect 495360 2922 495388 9114
rect 495544 3194 495572 9250
rect 496464 3534 496492 9522
rect 497476 9178 497504 12022
rect 497464 9172 497516 9178
rect 497464 9114 497516 9120
rect 496912 9104 496964 9110
rect 496912 9046 496964 9052
rect 496452 3528 496504 3534
rect 496452 3470 496504 3476
rect 495532 3188 495584 3194
rect 495532 3130 495584 3136
rect 496924 3058 496952 9046
rect 498200 8696 498252 8702
rect 498200 8638 498252 8644
rect 498212 4010 498240 8638
rect 498580 8566 498608 12022
rect 499500 9586 499528 12022
rect 499488 9580 499540 9586
rect 499488 9522 499540 9528
rect 499672 9512 499724 9518
rect 499672 9454 499724 9460
rect 498568 8560 498620 8566
rect 498568 8502 498620 8508
rect 498200 4004 498252 4010
rect 498200 3946 498252 3952
rect 499684 3534 499712 9454
rect 500788 9110 500816 12022
rect 501892 9654 501920 12022
rect 501880 9648 501932 9654
rect 501880 9590 501932 9596
rect 502996 9518 503024 12022
rect 502984 9512 503036 9518
rect 502984 9454 503036 9460
rect 503628 9444 503680 9450
rect 503628 9386 503680 9392
rect 500776 9104 500828 9110
rect 500776 9046 500828 9052
rect 500960 8968 501012 8974
rect 500960 8910 501012 8916
rect 499396 3528 499448 3534
rect 499396 3470 499448 3476
rect 499672 3528 499724 3534
rect 499672 3470 499724 3476
rect 498200 3188 498252 3194
rect 498200 3130 498252 3136
rect 495900 3052 495952 3058
rect 495900 2994 495952 3000
rect 496912 3052 496964 3058
rect 496912 2994 496964 3000
rect 495348 2916 495400 2922
rect 495348 2858 495400 2864
rect 495912 480 495940 2994
rect 497096 2916 497148 2922
rect 497096 2858 497148 2864
rect 497108 480 497136 2858
rect 498212 480 498240 3130
rect 499408 480 499436 3470
rect 500972 3330 501000 8910
rect 501052 8900 501104 8906
rect 501052 8842 501104 8848
rect 501064 3466 501092 8842
rect 501788 4004 501840 4010
rect 501788 3946 501840 3952
rect 501052 3460 501104 3466
rect 501052 3402 501104 3408
rect 500960 3324 501012 3330
rect 500960 3266 501012 3272
rect 500592 3052 500644 3058
rect 500592 2994 500644 3000
rect 500604 480 500632 2994
rect 501800 480 501828 3946
rect 502984 3528 503036 3534
rect 502984 3470 503036 3476
rect 502996 480 503024 3470
rect 503640 3262 503668 9386
rect 504100 9314 504128 12022
rect 505020 9450 505048 12022
rect 505008 9444 505060 9450
rect 505008 9386 505060 9392
rect 504088 9308 504140 9314
rect 504088 9250 504140 9256
rect 505008 9240 505060 9246
rect 505008 9182 505060 9188
rect 504180 3324 504232 3330
rect 504180 3266 504232 3272
rect 503628 3256 503680 3262
rect 503628 3198 503680 3204
rect 504192 480 504220 3266
rect 505020 3194 505048 9182
rect 506308 8906 506336 12022
rect 507412 9246 507440 12022
rect 507400 9240 507452 9246
rect 507400 9182 507452 9188
rect 506480 9036 506532 9042
rect 506480 8978 506532 8984
rect 506296 8900 506348 8906
rect 506296 8842 506348 8848
rect 505560 8628 505612 8634
rect 505560 8570 505612 8576
rect 505572 3534 505600 8570
rect 505560 3528 505612 3534
rect 505560 3470 505612 3476
rect 506492 3466 506520 8978
rect 508516 8838 508544 12022
rect 508504 8832 508556 8838
rect 508504 8774 508556 8780
rect 507860 8764 507912 8770
rect 507860 8706 507912 8712
rect 506756 8492 506808 8498
rect 506756 8434 506808 8440
rect 506768 4146 506796 8434
rect 506756 4140 506808 4146
rect 506756 4082 506808 4088
rect 507872 3602 507900 8706
rect 509620 8498 509648 12022
rect 510160 9376 510212 9382
rect 510160 9318 510212 9324
rect 509608 8492 509660 8498
rect 509608 8434 509660 8440
rect 507860 3596 507912 3602
rect 507860 3538 507912 3544
rect 508872 3528 508924 3534
rect 508872 3470 508924 3476
rect 505376 3460 505428 3466
rect 505376 3402 505428 3408
rect 506480 3460 506532 3466
rect 506480 3402 506532 3408
rect 505008 3188 505060 3194
rect 505008 3130 505060 3136
rect 505388 480 505416 3402
rect 506480 3256 506532 3262
rect 506480 3198 506532 3204
rect 506492 480 506520 3198
rect 507676 3188 507728 3194
rect 507676 3130 507728 3136
rect 507688 480 507716 3130
rect 508884 480 508912 3470
rect 510068 3460 510120 3466
rect 510068 3402 510120 3408
rect 510080 480 510108 3402
rect 510172 3330 510200 9318
rect 510540 8974 510568 12022
rect 510712 9172 510764 9178
rect 510712 9114 510764 9120
rect 510528 8968 510580 8974
rect 510528 8910 510580 8916
rect 510724 3466 510752 9114
rect 511828 8770 511856 12022
rect 511816 8764 511868 8770
rect 511816 8706 511868 8712
rect 512932 8702 512960 12022
rect 513196 9580 513248 9586
rect 513196 9522 513248 9528
rect 512920 8696 512972 8702
rect 512920 8638 512972 8644
rect 511264 4140 511316 4146
rect 511264 4082 511316 4088
rect 510712 3460 510764 3466
rect 510712 3402 510764 3408
rect 510160 3324 510212 3330
rect 510160 3266 510212 3272
rect 511276 480 511304 4082
rect 512460 3596 512512 3602
rect 512460 3538 512512 3544
rect 512472 480 512500 3538
rect 513208 3398 513236 9522
rect 514036 9382 514064 12022
rect 514024 9376 514076 9382
rect 514024 9318 514076 9324
rect 514668 9104 514720 9110
rect 514668 9046 514720 9052
rect 513288 8560 513340 8566
rect 513288 8502 513340 8508
rect 513300 3534 513328 8502
rect 513288 3528 513340 3534
rect 513288 3470 513340 3476
rect 513196 3392 513248 3398
rect 513196 3334 513248 3340
rect 513564 3324 513616 3330
rect 513564 3266 513616 3272
rect 513576 480 513604 3266
rect 514680 3194 514708 9046
rect 515140 8634 515168 12022
rect 515956 9648 516008 9654
rect 515956 9590 516008 9596
rect 515128 8628 515180 8634
rect 515128 8570 515180 8576
rect 515968 6914 515996 9590
rect 516060 9586 516088 12022
rect 516048 9580 516100 9586
rect 516048 9522 516100 9528
rect 516508 9512 516560 9518
rect 516508 9454 516560 9460
rect 515968 6886 516088 6914
rect 516060 3602 516088 6886
rect 516520 4146 516548 9454
rect 517348 9178 517376 12022
rect 518452 9654 518480 12022
rect 518440 9648 518492 9654
rect 518440 9590 518492 9596
rect 517612 9444 517664 9450
rect 517612 9386 517664 9392
rect 517520 9308 517572 9314
rect 517520 9250 517572 9256
rect 517336 9172 517388 9178
rect 517336 9114 517388 9120
rect 516508 4140 516560 4146
rect 516508 4082 516560 4088
rect 516048 3596 516100 3602
rect 516048 3538 516100 3544
rect 517532 3534 517560 9250
rect 515956 3528 516008 3534
rect 515956 3470 516008 3476
rect 517520 3528 517572 3534
rect 517520 3470 517572 3476
rect 514760 3460 514812 3466
rect 514760 3402 514812 3408
rect 514668 3188 514720 3194
rect 514668 3130 514720 3136
rect 514772 480 514800 3402
rect 515968 480 515996 3470
rect 517624 3466 517652 9386
rect 519556 9314 519584 12022
rect 519544 9308 519596 9314
rect 519544 9250 519596 9256
rect 520464 9240 520516 9246
rect 520464 9182 520516 9188
rect 518900 8900 518952 8906
rect 518900 8842 518952 8848
rect 517612 3460 517664 3466
rect 517612 3402 517664 3408
rect 517152 3392 517204 3398
rect 517152 3334 517204 3340
rect 517164 480 517192 3334
rect 518912 3262 518940 8842
rect 519544 3596 519596 3602
rect 519544 3538 519596 3544
rect 518900 3256 518952 3262
rect 518900 3198 518952 3204
rect 518348 3188 518400 3194
rect 518348 3130 518400 3136
rect 518360 480 518388 3130
rect 519556 480 519584 3538
rect 520476 3398 520504 9182
rect 520660 9042 520688 12022
rect 520648 9036 520700 9042
rect 520648 8978 520700 8984
rect 521580 8906 521608 12022
rect 522868 9450 522896 12022
rect 522856 9444 522908 9450
rect 522856 9386 522908 9392
rect 523972 9110 524000 12022
rect 525076 9246 525104 12022
rect 525812 12022 525872 12050
rect 525996 12022 526976 12050
rect 528080 12022 528324 12050
rect 529184 12022 529520 12050
rect 530288 12022 530624 12050
rect 531392 12022 531544 12050
rect 525064 9240 525116 9246
rect 525064 9182 525116 9188
rect 523960 9104 524012 9110
rect 523960 9046 524012 9052
rect 524236 8968 524288 8974
rect 524236 8910 524288 8916
rect 521568 8900 521620 8906
rect 521568 8842 521620 8848
rect 522948 8832 523000 8838
rect 522948 8774 523000 8780
rect 520740 4140 520792 4146
rect 520740 4082 520792 4088
rect 520464 3392 520516 3398
rect 520464 3334 520516 3340
rect 520752 480 520780 4082
rect 521844 3528 521896 3534
rect 521844 3470 521896 3476
rect 521856 480 521884 3470
rect 522960 3194 522988 8774
rect 524248 4078 524276 8910
rect 525812 8770 525840 12022
rect 525708 8764 525760 8770
rect 525708 8706 525760 8712
rect 525800 8764 525852 8770
rect 525800 8706 525852 8712
rect 524328 8492 524380 8498
rect 524328 8434 524380 8440
rect 524236 4072 524288 4078
rect 524236 4014 524288 4020
rect 524340 3534 524368 8434
rect 525720 4146 525748 8706
rect 525708 4140 525760 4146
rect 525708 4082 525760 4088
rect 524328 3528 524380 3534
rect 524328 3470 524380 3476
rect 523040 3460 523092 3466
rect 523040 3402 523092 3408
rect 522948 3188 523000 3194
rect 522948 3130 523000 3136
rect 523052 480 523080 3402
rect 525432 3392 525484 3398
rect 525996 3369 526024 12022
rect 528296 9518 528324 12022
rect 528652 9580 528704 9586
rect 528652 9522 528704 9528
rect 528284 9512 528336 9518
rect 528284 9454 528336 9460
rect 527916 9376 527968 9382
rect 527916 9318 527968 9324
rect 526444 8696 526496 8702
rect 526444 8638 526496 8644
rect 526456 3602 526484 8638
rect 527928 3738 527956 9318
rect 528560 8628 528612 8634
rect 528560 8570 528612 8576
rect 527916 3732 527968 3738
rect 527916 3674 527968 3680
rect 526444 3596 526496 3602
rect 526444 3538 526496 3544
rect 528572 3534 528600 8570
rect 527824 3528 527876 3534
rect 527824 3470 527876 3476
rect 528560 3528 528612 3534
rect 528560 3470 528612 3476
rect 525432 3334 525484 3340
rect 525982 3360 526038 3369
rect 524236 3256 524288 3262
rect 524236 3198 524288 3204
rect 524248 480 524276 3198
rect 525444 480 525472 3334
rect 525982 3295 526038 3304
rect 526628 3188 526680 3194
rect 526628 3130 526680 3136
rect 526640 480 526668 3130
rect 527836 480 527864 3470
rect 528664 2922 528692 9522
rect 529492 9382 529520 12022
rect 529480 9376 529532 9382
rect 529480 9318 529532 9324
rect 530032 9172 530084 9178
rect 530032 9114 530084 9120
rect 529020 4072 529072 4078
rect 529020 4014 529072 4020
rect 528652 2916 528704 2922
rect 528652 2858 528704 2864
rect 529032 480 529060 4014
rect 530044 3398 530072 9114
rect 530596 8974 530624 12022
rect 530584 8968 530636 8974
rect 530584 8910 530636 8916
rect 531516 8838 531544 12022
rect 531608 12022 532496 12050
rect 532804 12022 533600 12050
rect 534704 12022 535040 12050
rect 535808 12022 536144 12050
rect 536912 12022 537248 12050
rect 538016 12022 538168 12050
rect 539120 12022 539456 12050
rect 540224 12022 540560 12050
rect 541328 12022 541664 12050
rect 542432 12022 542768 12050
rect 543536 12022 543688 12050
rect 544640 12022 544976 12050
rect 531504 8832 531556 8838
rect 531504 8774 531556 8780
rect 531608 6914 531636 12022
rect 532608 9648 532660 9654
rect 532608 9590 532660 9596
rect 531424 6886 531636 6914
rect 530124 4140 530176 4146
rect 530124 4082 530176 4088
rect 530032 3392 530084 3398
rect 530032 3334 530084 3340
rect 530136 480 530164 4082
rect 531424 3602 531452 6886
rect 532516 3732 532568 3738
rect 532516 3674 532568 3680
rect 531320 3596 531372 3602
rect 531320 3538 531372 3544
rect 531412 3596 531464 3602
rect 531412 3538 531464 3544
rect 531332 480 531360 3538
rect 532528 480 532556 3674
rect 532620 3466 532648 9590
rect 532804 3777 532832 12022
rect 535012 9586 535040 12022
rect 535000 9580 535052 9586
rect 535000 9522 535052 9528
rect 536012 9444 536064 9450
rect 536012 9386 536064 9392
rect 533988 9308 534040 9314
rect 533988 9250 534040 9256
rect 534000 4010 534028 9250
rect 534908 9036 534960 9042
rect 534908 8978 534960 8984
rect 533988 4004 534040 4010
rect 533988 3946 534040 3952
rect 534920 3942 534948 8978
rect 535368 8900 535420 8906
rect 535368 8842 535420 8848
rect 535380 4146 535408 8842
rect 535368 4140 535420 4146
rect 535368 4082 535420 4088
rect 534908 3936 534960 3942
rect 534908 3878 534960 3884
rect 536024 3874 536052 9386
rect 536116 3913 536144 12022
rect 537220 9042 537248 12022
rect 538140 9314 538168 12022
rect 538128 9308 538180 9314
rect 538128 9250 538180 9256
rect 538864 9240 538916 9246
rect 538864 9182 538916 9188
rect 538036 9104 538088 9110
rect 538036 9046 538088 9052
rect 537208 9036 537260 9042
rect 537208 8978 537260 8984
rect 536102 3904 536158 3913
rect 536012 3868 536064 3874
rect 536102 3839 536158 3848
rect 536012 3810 536064 3816
rect 538048 3806 538076 9046
rect 538404 4004 538456 4010
rect 538404 3946 538456 3952
rect 538036 3800 538088 3806
rect 532790 3768 532846 3777
rect 538036 3742 538088 3748
rect 532790 3703 532846 3712
rect 533712 3528 533764 3534
rect 533712 3470 533764 3476
rect 532608 3460 532660 3466
rect 532608 3402 532660 3408
rect 533724 480 533752 3470
rect 537208 3460 537260 3466
rect 537208 3402 537260 3408
rect 536104 3392 536156 3398
rect 536104 3334 536156 3340
rect 534908 2916 534960 2922
rect 534908 2858 534960 2864
rect 534920 480 534948 2858
rect 536116 480 536144 3334
rect 537220 480 537248 3402
rect 538416 480 538444 3946
rect 538876 3602 538904 9182
rect 539428 4078 539456 12022
rect 539692 8764 539744 8770
rect 539692 8706 539744 8712
rect 539416 4072 539468 4078
rect 539416 4014 539468 4020
rect 539600 3936 539652 3942
rect 539600 3878 539652 3884
rect 538864 3596 538916 3602
rect 538864 3538 538916 3544
rect 539612 480 539640 3878
rect 539704 2990 539732 8706
rect 540532 4010 540560 12022
rect 540980 9512 541032 9518
rect 540980 9454 541032 9460
rect 540796 4140 540848 4146
rect 540796 4082 540848 4088
rect 540520 4004 540572 4010
rect 540520 3946 540572 3952
rect 539692 2984 539744 2990
rect 539692 2926 539744 2932
rect 540808 480 540836 4082
rect 540992 3262 541020 9454
rect 541636 9178 541664 12022
rect 542360 9376 542412 9382
rect 542360 9318 542412 9324
rect 541624 9172 541676 9178
rect 541624 9114 541676 9120
rect 542372 3874 542400 9318
rect 542740 4146 542768 12022
rect 542728 4140 542780 4146
rect 542728 4082 542780 4088
rect 541992 3868 542044 3874
rect 541992 3810 542044 3816
rect 542360 3868 542412 3874
rect 542360 3810 542412 3816
rect 540980 3256 541032 3262
rect 540980 3198 541032 3204
rect 542004 480 542032 3810
rect 543188 3800 543240 3806
rect 543188 3742 543240 3748
rect 543200 480 543228 3742
rect 543660 3641 543688 12022
rect 544948 9110 544976 12022
rect 545132 12022 545744 12050
rect 546512 12022 546848 12050
rect 544936 9104 544988 9110
rect 544936 9046 544988 9052
rect 545028 8968 545080 8974
rect 545028 8910 545080 8916
rect 545040 3942 545068 8910
rect 545028 3936 545080 3942
rect 545028 3878 545080 3884
rect 543646 3632 543702 3641
rect 543646 3567 543702 3576
rect 544384 3596 544436 3602
rect 544384 3538 544436 3544
rect 544396 480 544424 3538
rect 545132 3398 545160 12022
rect 545764 8832 545816 8838
rect 545764 8774 545816 8780
rect 545776 3738 545804 8774
rect 546512 4049 546540 12022
rect 547938 11778 547966 12036
rect 548076 12022 549056 12050
rect 549364 12022 550160 12050
rect 550652 12022 551264 12050
rect 552032 12022 552368 12050
rect 553412 12022 553472 12050
rect 553688 12022 554576 12050
rect 554792 12022 555680 12050
rect 556172 12022 556784 12050
rect 557552 12022 557888 12050
rect 558932 12022 558992 12050
rect 559300 12022 560096 12050
rect 560312 12022 561200 12050
rect 547938 11750 548012 11778
rect 547880 9580 547932 9586
rect 547880 9522 547932 9528
rect 546498 4040 546554 4049
rect 546498 3975 546554 3984
rect 545764 3732 545816 3738
rect 545764 3674 545816 3680
rect 547892 3602 547920 9522
rect 547984 8974 548012 11750
rect 547972 8968 548024 8974
rect 547972 8910 548024 8916
rect 547880 3596 547932 3602
rect 547880 3538 547932 3544
rect 545120 3392 545172 3398
rect 548076 3369 548104 12022
rect 549076 3868 549128 3874
rect 549076 3810 549128 3816
rect 545120 3334 545172 3340
rect 546682 3360 546738 3369
rect 546682 3295 546738 3304
rect 548062 3360 548118 3369
rect 548062 3295 548118 3304
rect 545488 2984 545540 2990
rect 545488 2926 545540 2932
rect 545500 480 545528 2926
rect 546696 480 546724 3295
rect 547880 3256 547932 3262
rect 547880 3198 547932 3204
rect 547892 480 547920 3198
rect 549088 480 549116 3810
rect 549364 3505 549392 12022
rect 550272 3936 550324 3942
rect 550272 3878 550324 3884
rect 549350 3496 549406 3505
rect 549350 3431 549406 3440
rect 550284 480 550312 3878
rect 550652 3806 550680 12022
rect 551836 9308 551888 9314
rect 551836 9250 551888 9256
rect 550640 3800 550692 3806
rect 550640 3742 550692 3748
rect 551468 3732 551520 3738
rect 551468 3674 551520 3680
rect 551480 480 551508 3674
rect 551848 3670 551876 9250
rect 551928 9036 551980 9042
rect 551928 8978 551980 8984
rect 551836 3664 551888 3670
rect 551836 3606 551888 3612
rect 551940 3534 551968 8978
rect 552032 3942 552060 12022
rect 553412 3942 553440 12022
rect 553688 6914 553716 12022
rect 553504 6886 553716 6914
rect 552020 3936 552072 3942
rect 552020 3878 552072 3884
rect 553216 3936 553268 3942
rect 553216 3878 553268 3884
rect 553400 3936 553452 3942
rect 553400 3878 553452 3884
rect 552756 3800 552808 3806
rect 552756 3742 552808 3748
rect 551928 3528 551980 3534
rect 551928 3470 551980 3476
rect 552768 3466 552796 3742
rect 552664 3460 552716 3466
rect 552664 3402 552716 3408
rect 552756 3460 552808 3466
rect 552756 3402 552808 3408
rect 552676 480 552704 3402
rect 553228 3330 553256 3878
rect 553504 3874 553532 6886
rect 553492 3868 553544 3874
rect 553492 3810 553544 3816
rect 554792 3806 554820 12022
rect 555424 9172 555476 9178
rect 555424 9114 555476 9120
rect 554780 3800 554832 3806
rect 553766 3768 553822 3777
rect 554780 3742 554832 3748
rect 553766 3703 553822 3712
rect 553216 3324 553268 3330
rect 553216 3266 553268 3272
rect 553780 480 553808 3703
rect 554964 3596 555016 3602
rect 554964 3538 555016 3544
rect 554976 480 555004 3538
rect 555436 3194 555464 9114
rect 556172 3738 556200 12022
rect 556342 3904 556398 3913
rect 556342 3839 556398 3848
rect 556160 3732 556212 3738
rect 556160 3674 556212 3680
rect 555424 3188 555476 3194
rect 555424 3130 555476 3136
rect 479310 354 479422 480
rect 478892 326 479422 354
rect 479310 -960 479422 326
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 218 556242 480
rect 556356 218 556384 3839
rect 557356 3528 557408 3534
rect 557356 3470 557408 3476
rect 557368 480 557396 3470
rect 557552 3466 557580 12022
rect 557632 9104 557684 9110
rect 557632 9046 557684 9052
rect 557540 3460 557592 3466
rect 557540 3402 557592 3408
rect 557644 3398 557672 9046
rect 558552 3664 558604 3670
rect 558552 3606 558604 3612
rect 557632 3392 557684 3398
rect 557632 3334 557684 3340
rect 558564 480 558592 3606
rect 558932 3602 558960 12022
rect 559300 6914 559328 12022
rect 559024 6886 559328 6914
rect 559024 3777 559052 6886
rect 559748 4072 559800 4078
rect 559748 4014 559800 4020
rect 559010 3768 559066 3777
rect 559010 3703 559066 3712
rect 558920 3596 558972 3602
rect 558920 3538 558972 3544
rect 559760 480 559788 4014
rect 560312 3670 560340 12022
rect 568488 8968 568540 8974
rect 568488 8910 568540 8916
rect 563244 4140 563296 4146
rect 563244 4082 563296 4088
rect 560852 4004 560904 4010
rect 560852 3946 560904 3952
rect 560300 3664 560352 3670
rect 560300 3606 560352 3612
rect 560864 480 560892 3946
rect 562048 3188 562100 3194
rect 562048 3130 562100 3136
rect 562060 480 562088 3130
rect 563256 480 563284 4082
rect 568026 4040 568082 4049
rect 568026 3975 568082 3984
rect 564438 3632 564494 3641
rect 564438 3567 564494 3576
rect 564452 480 564480 3567
rect 565636 3392 565688 3398
rect 565636 3334 565688 3340
rect 565648 480 565676 3334
rect 566832 3256 566884 3262
rect 566832 3198 566884 3204
rect 566844 480 566872 3198
rect 568040 480 568068 3975
rect 568500 2802 568528 8910
rect 578896 6633 578924 19314
rect 578882 6624 578938 6633
rect 578882 6559 578938 6568
rect 575112 3936 575164 3942
rect 575112 3878 575164 3884
rect 572720 3528 572772 3534
rect 571522 3496 571578 3505
rect 572720 3470 572772 3476
rect 571522 3431 571578 3440
rect 570326 3360 570382 3369
rect 570326 3295 570382 3304
rect 568500 2774 568712 2802
rect 556130 190 556384 218
rect 556130 -960 556242 190
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 568684 354 568712 2774
rect 570340 480 570368 3295
rect 571536 480 571564 3431
rect 572732 480 572760 3470
rect 573916 3324 573968 3330
rect 573916 3266 573968 3272
rect 573928 480 573956 3266
rect 575124 480 575152 3878
rect 576308 3868 576360 3874
rect 576308 3810 576360 3816
rect 576320 480 576348 3810
rect 577412 3800 577464 3806
rect 577412 3742 577464 3748
rect 582194 3768 582250 3777
rect 577424 480 577452 3742
rect 578608 3732 578660 3738
rect 582194 3703 582250 3712
rect 578608 3674 578660 3680
rect 578620 480 578648 3674
rect 581000 3596 581052 3602
rect 581000 3538 581052 3544
rect 579804 3460 579856 3466
rect 579804 3402 579856 3408
rect 579816 480 579844 3402
rect 581012 480 581040 3538
rect 582208 480 582236 3703
rect 583392 3664 583444 3670
rect 583392 3606 583444 3612
rect 583404 480 583432 3606
rect 569102 354 569214 480
rect 568684 326 569214 354
rect 569102 -960 569214 326
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3422 697312 3478 697368
rect 3514 684256 3570 684312
rect 580170 697176 580226 697232
rect 3606 671200 3662 671256
rect 3422 658144 3478 658200
rect 580170 683848 580226 683904
rect 569222 670520 569278 670576
rect 9402 669568 9458 669624
rect 580170 670692 580172 670712
rect 580172 670692 580224 670712
rect 580224 670692 580226 670712
rect 569314 658008 569370 658064
rect 9402 657328 9458 657384
rect 3514 645088 3570 645144
rect 9402 645088 9458 645144
rect 580170 670656 580226 670692
rect 580170 657328 580226 657384
rect 569406 645496 569462 645552
rect 580170 644000 580226 644056
rect 569222 632984 569278 633040
rect 8666 632848 8722 632904
rect 3606 632032 3662 632088
rect 3422 619112 3478 619168
rect 8666 620608 8722 620664
rect 9402 608368 9458 608424
rect 580170 630808 580226 630864
rect 569314 620472 569370 620528
rect 580170 617480 580226 617536
rect 569222 607960 569278 608016
rect 3514 606056 3570 606112
rect 2778 593000 2834 593056
rect 9402 596148 9458 596184
rect 9402 596128 9404 596148
rect 9404 596128 9456 596148
rect 9456 596128 9458 596148
rect 580170 604152 580226 604208
rect 569314 595448 569370 595504
rect 2962 579944 3018 580000
rect 3422 566888 3478 566944
rect 9402 583888 9458 583944
rect 8850 571648 8906 571704
rect 579802 590960 579858 591016
rect 569406 582936 569462 582992
rect 580170 577632 580226 577688
rect 569222 570424 569278 570480
rect 9402 559408 9458 559464
rect 3514 553832 3570 553888
rect 3422 540776 3478 540832
rect 9402 547168 9458 547224
rect 579802 564304 579858 564360
rect 569314 557912 569370 557968
rect 580170 551112 580226 551168
rect 569222 545400 569278 545456
rect 3422 527856 3478 527912
rect 3422 514820 3478 514856
rect 3422 514800 3424 514820
rect 3424 514800 3476 514820
rect 3476 514800 3478 514820
rect 9402 534928 9458 534984
rect 7654 522688 7710 522744
rect 580170 537784 580226 537840
rect 569314 532888 569370 532944
rect 580170 524476 580226 524512
rect 580170 524456 580172 524476
rect 580172 524456 580224 524476
rect 580224 524456 580226 524476
rect 569222 520376 569278 520432
rect 7562 510448 7618 510504
rect 3054 501744 3110 501800
rect 8942 498208 8998 498264
rect 3422 488708 3478 488744
rect 3422 488688 3424 488708
rect 3424 488688 3476 488708
rect 3476 488688 3478 488708
rect 3422 475652 3478 475688
rect 3422 475632 3424 475652
rect 3424 475632 3476 475652
rect 3476 475632 3478 475652
rect 580170 511264 580226 511320
rect 569314 507864 569370 507920
rect 579894 497936 579950 497992
rect 569222 495352 569278 495408
rect 9034 485968 9090 486024
rect 580630 484608 580686 484664
rect 569866 482840 569922 482896
rect 8942 473728 8998 473784
rect 3422 462596 3478 462632
rect 3422 462576 3424 462596
rect 3424 462576 3476 462596
rect 3476 462576 3478 462596
rect 2778 449520 2834 449576
rect 569866 470328 569922 470384
rect 9034 461488 9090 461544
rect 579986 471416 580042 471472
rect 580262 458088 580318 458144
rect 569866 457852 569868 457872
rect 569868 457852 569920 457872
rect 569920 457852 569922 457872
rect 569866 457816 569922 457852
rect 8942 449248 8998 449304
rect 569130 445304 569186 445360
rect 580354 444760 580410 444816
rect 9402 437008 9458 437064
rect 2962 436600 3018 436656
rect 569314 432792 569370 432848
rect 580170 431568 580226 431624
rect 9402 424768 9458 424824
rect 3422 423544 3478 423600
rect 569222 420280 569278 420336
rect 580170 418240 580226 418296
rect 7562 412528 7618 412584
rect 3146 410488 3202 410544
rect 569222 407768 569278 407824
rect 580170 404912 580226 404968
rect 7562 400288 7618 400344
rect 3422 397468 3424 397488
rect 3424 397468 3476 397488
rect 3476 397468 3478 397488
rect 3422 397432 3478 397468
rect 569130 395256 569186 395312
rect 578882 391720 578938 391776
rect 7562 388048 7618 388104
rect 3422 384376 3478 384432
rect 569866 382744 569922 382800
rect 578882 378392 578938 378448
rect 7562 375808 7618 375864
rect 3422 371340 3478 371376
rect 3422 371320 3424 371340
rect 3424 371320 3476 371340
rect 3476 371320 3478 371340
rect 569590 370232 569646 370288
rect 579618 365064 579674 365120
rect 7562 363568 7618 363624
rect 2778 358400 2834 358456
rect 569682 357720 569738 357776
rect 579526 351872 579582 351928
rect 8666 351328 8722 351384
rect 4066 345344 4122 345400
rect 569682 345208 569738 345264
rect 9402 339088 9458 339144
rect 580170 338544 580226 338600
rect 569222 332696 569278 332752
rect 3054 332288 3110 332344
rect 9402 326848 9458 326904
rect 580170 325216 580226 325272
rect 568670 320184 568726 320240
rect 3422 319232 3478 319288
rect 9402 314628 9458 314664
rect 9402 314608 9404 314628
rect 9404 314608 9456 314628
rect 9456 314608 9458 314628
rect 580170 312024 580226 312080
rect 568946 307672 569002 307728
rect 3422 306196 3478 306232
rect 3422 306176 3424 306196
rect 3424 306176 3476 306196
rect 3476 306176 3478 306196
rect 9402 302368 9458 302424
rect 580354 298696 580410 298752
rect 569866 295160 569922 295216
rect 3422 293120 3478 293176
rect 9402 290128 9458 290184
rect 580170 285368 580226 285424
rect 569866 282684 569868 282704
rect 569868 282684 569920 282704
rect 569920 282684 569922 282704
rect 569866 282648 569922 282684
rect 3422 280064 3478 280120
rect 9218 277888 9274 277944
rect 579802 272176 579858 272232
rect 569314 270172 569316 270192
rect 569316 270172 569368 270192
rect 569368 270172 569370 270192
rect 569314 270136 569370 270172
rect 3054 267144 3110 267200
rect 9402 265648 9458 265704
rect 579710 258848 579766 258904
rect 569130 257624 569186 257680
rect 3422 254108 3478 254144
rect 3422 254088 3424 254108
rect 3424 254088 3476 254108
rect 3476 254088 3478 254108
rect 9402 253408 9458 253464
rect 580170 245520 580226 245576
rect 568670 245112 568726 245168
rect 9402 241168 9458 241224
rect 3422 241032 3478 241088
rect 569866 232600 569922 232656
rect 580170 232328 580226 232384
rect 8850 228928 8906 228984
rect 3422 227996 3478 228032
rect 3422 227976 3424 227996
rect 3424 227976 3476 227996
rect 3476 227976 3478 227996
rect 569498 220088 569554 220144
rect 580446 219000 580502 219056
rect 8206 216688 8262 216744
rect 3422 214956 3424 214976
rect 3424 214956 3476 214976
rect 3476 214956 3478 214976
rect 3422 214920 3478 214956
rect 569866 207576 569922 207632
rect 579526 205672 579582 205728
rect 8206 204448 8262 204504
rect 3330 201864 3386 201920
rect 569314 195064 569370 195120
rect 579526 192480 579582 192536
rect 8206 192208 8262 192264
rect 3422 188844 3424 188864
rect 3424 188844 3476 188864
rect 3476 188844 3478 188864
rect 3422 188808 3478 188844
rect 569406 182552 569462 182608
rect 8206 179968 8262 180024
rect 580262 179152 580318 179208
rect 3422 175888 3478 175944
rect 569866 170040 569922 170096
rect 8206 167728 8262 167784
rect 579986 165824 580042 165880
rect 3514 162832 3570 162888
rect 569866 157528 569922 157584
rect 8942 155488 8998 155544
rect 579526 152632 579582 152688
rect 3422 149776 3478 149832
rect 569866 145016 569922 145072
rect 8298 143248 8354 143304
rect 578882 139304 578938 139360
rect 3238 136720 3294 136776
rect 569866 132524 569922 132560
rect 569866 132504 569868 132524
rect 569868 132504 569920 132524
rect 569920 132504 569922 132524
rect 9034 131008 9090 131064
rect 4066 123664 4122 123720
rect 579618 125976 579674 126032
rect 568670 119992 568726 120048
rect 9402 118768 9458 118824
rect 578882 112784 578938 112840
rect 2778 110608 2834 110664
rect 569682 107480 569738 107536
rect 9402 106528 9458 106584
rect 578882 99456 578938 99512
rect 2778 97552 2834 97608
rect 569682 94968 569738 95024
rect 9402 94288 9458 94344
rect 580170 86128 580226 86184
rect 2778 84632 2834 84688
rect 569682 82456 569738 82512
rect 8942 82048 8998 82104
rect 578882 72936 578938 72992
rect 3422 71612 3424 71632
rect 3424 71612 3476 71632
rect 3476 71612 3478 71632
rect 3422 71576 3478 71612
rect 569590 69944 569646 70000
rect 8942 69808 8998 69864
rect 578882 59608 578938 59664
rect 3146 58520 3202 58576
rect 8850 57568 8906 57624
rect 569130 57432 569186 57488
rect 580170 46280 580226 46336
rect 2778 45500 2780 45520
rect 2780 45500 2832 45520
rect 2832 45500 2834 45520
rect 2778 45464 2834 45500
rect 9402 45328 9458 45384
rect 569866 44920 569922 44976
rect 9034 33088 9090 33144
rect 578882 33088 578938 33144
rect 2778 32408 2834 32464
rect 569498 32408 569554 32464
rect 8942 20848 8998 20904
rect 2778 19352 2834 19408
rect 569866 19896 569922 19952
rect 578974 19760 579030 19816
rect 3422 6468 3424 6488
rect 3424 6468 3476 6488
rect 3476 6468 3478 6488
rect 3422 6432 3478 6468
rect 525982 3304 526038 3360
rect 536102 3848 536158 3904
rect 532790 3712 532846 3768
rect 543646 3576 543702 3632
rect 546498 3984 546554 4040
rect 546682 3304 546738 3360
rect 548062 3304 548118 3360
rect 549350 3440 549406 3496
rect 553766 3712 553822 3768
rect 556342 3848 556398 3904
rect 559010 3712 559066 3768
rect 568026 3984 568082 4040
rect 564438 3576 564494 3632
rect 578882 6568 578938 6624
rect 571522 3440 571578 3496
rect 570326 3304 570382 3360
rect 582194 3712 582250 3768
<< metal3 >>
rect -960 697370 480 697460
rect 3417 697370 3483 697373
rect -960 697368 3483 697370
rect -960 697312 3422 697368
rect 3478 697312 3483 697368
rect -960 697310 3483 697312
rect -960 697220 480 697310
rect 3417 697307 3483 697310
rect 580165 697234 580231 697237
rect 583520 697234 584960 697324
rect 580165 697232 584960 697234
rect 580165 697176 580170 697232
rect 580226 697176 584960 697232
rect 580165 697174 584960 697176
rect 580165 697171 580231 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 3509 684314 3575 684317
rect -960 684312 3575 684314
rect -960 684256 3514 684312
rect 3570 684256 3575 684312
rect -960 684254 3575 684256
rect -960 684164 480 684254
rect 3509 684251 3575 684254
rect 580165 683906 580231 683909
rect 583520 683906 584960 683996
rect 580165 683904 584960 683906
rect 580165 683848 580170 683904
rect 580226 683848 584960 683904
rect 580165 683846 584960 683848
rect 580165 683843 580231 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 3601 671258 3667 671261
rect -960 671256 3667 671258
rect -960 671200 3606 671256
rect 3662 671200 3667 671256
rect -960 671198 3667 671200
rect -960 671108 480 671198
rect 3601 671195 3667 671198
rect 580165 670714 580231 670717
rect 583520 670714 584960 670804
rect 580165 670712 584960 670714
rect 580165 670656 580170 670712
rect 580226 670656 584960 670712
rect 580165 670654 584960 670656
rect 580165 670651 580231 670654
rect 569217 670578 569283 670581
rect 566076 670576 569283 670578
rect 566076 670520 569222 670576
rect 569278 670520 569283 670576
rect 583520 670564 584960 670654
rect 566076 670518 569283 670520
rect 569217 670515 569283 670518
rect 9397 669626 9463 669629
rect 9397 669624 12052 669626
rect 9397 669568 9402 669624
rect 9458 669568 12052 669624
rect 9397 669566 12052 669568
rect 9397 669563 9463 669566
rect -960 658202 480 658292
rect 3417 658202 3483 658205
rect -960 658200 3483 658202
rect -960 658144 3422 658200
rect 3478 658144 3483 658200
rect -960 658142 3483 658144
rect -960 658052 480 658142
rect 3417 658139 3483 658142
rect 569309 658066 569375 658069
rect 566076 658064 569375 658066
rect 566076 658008 569314 658064
rect 569370 658008 569375 658064
rect 566076 658006 569375 658008
rect 569309 658003 569375 658006
rect 9397 657386 9463 657389
rect 580165 657386 580231 657389
rect 583520 657386 584960 657476
rect 9397 657384 12052 657386
rect 9397 657328 9402 657384
rect 9458 657328 12052 657384
rect 9397 657326 12052 657328
rect 580165 657384 584960 657386
rect 580165 657328 580170 657384
rect 580226 657328 584960 657384
rect 580165 657326 584960 657328
rect 9397 657323 9463 657326
rect 580165 657323 580231 657326
rect 583520 657236 584960 657326
rect 569401 645554 569467 645557
rect 566076 645552 569467 645554
rect 566076 645496 569406 645552
rect 569462 645496 569467 645552
rect 566076 645494 569467 645496
rect 569401 645491 569467 645494
rect -960 645146 480 645236
rect 3509 645146 3575 645149
rect -960 645144 3575 645146
rect -960 645088 3514 645144
rect 3570 645088 3575 645144
rect -960 645086 3575 645088
rect -960 644996 480 645086
rect 3509 645083 3575 645086
rect 9397 645146 9463 645149
rect 9397 645144 12052 645146
rect 9397 645088 9402 645144
rect 9458 645088 12052 645144
rect 9397 645086 12052 645088
rect 9397 645083 9463 645086
rect 580165 644058 580231 644061
rect 583520 644058 584960 644148
rect 580165 644056 584960 644058
rect 580165 644000 580170 644056
rect 580226 644000 584960 644056
rect 580165 643998 584960 644000
rect 580165 643995 580231 643998
rect 583520 643908 584960 643998
rect 569217 633042 569283 633045
rect 566076 633040 569283 633042
rect 566076 632984 569222 633040
rect 569278 632984 569283 633040
rect 566076 632982 569283 632984
rect 569217 632979 569283 632982
rect 8661 632906 8727 632909
rect 8661 632904 12052 632906
rect 8661 632848 8666 632904
rect 8722 632848 12052 632904
rect 8661 632846 12052 632848
rect 8661 632843 8727 632846
rect -960 632090 480 632180
rect 3601 632090 3667 632093
rect -960 632088 3667 632090
rect -960 632032 3606 632088
rect 3662 632032 3667 632088
rect -960 632030 3667 632032
rect -960 631940 480 632030
rect 3601 632027 3667 632030
rect 580165 630866 580231 630869
rect 583520 630866 584960 630956
rect 580165 630864 584960 630866
rect 580165 630808 580170 630864
rect 580226 630808 584960 630864
rect 580165 630806 584960 630808
rect 580165 630803 580231 630806
rect 583520 630716 584960 630806
rect 8661 620666 8727 620669
rect 8661 620664 12052 620666
rect 8661 620608 8666 620664
rect 8722 620608 12052 620664
rect 8661 620606 12052 620608
rect 8661 620603 8727 620606
rect 569309 620530 569375 620533
rect 566076 620528 569375 620530
rect 566076 620472 569314 620528
rect 569370 620472 569375 620528
rect 566076 620470 569375 620472
rect 569309 620467 569375 620470
rect -960 619170 480 619260
rect 3417 619170 3483 619173
rect -960 619168 3483 619170
rect -960 619112 3422 619168
rect 3478 619112 3483 619168
rect -960 619110 3483 619112
rect -960 619020 480 619110
rect 3417 619107 3483 619110
rect 580165 617538 580231 617541
rect 583520 617538 584960 617628
rect 580165 617536 584960 617538
rect 580165 617480 580170 617536
rect 580226 617480 584960 617536
rect 580165 617478 584960 617480
rect 580165 617475 580231 617478
rect 583520 617388 584960 617478
rect 9397 608426 9463 608429
rect 9397 608424 12052 608426
rect 9397 608368 9402 608424
rect 9458 608368 12052 608424
rect 9397 608366 12052 608368
rect 9397 608363 9463 608366
rect 569217 608018 569283 608021
rect 566076 608016 569283 608018
rect 566076 607960 569222 608016
rect 569278 607960 569283 608016
rect 566076 607958 569283 607960
rect 569217 607955 569283 607958
rect -960 606114 480 606204
rect 3509 606114 3575 606117
rect -960 606112 3575 606114
rect -960 606056 3514 606112
rect 3570 606056 3575 606112
rect -960 606054 3575 606056
rect -960 605964 480 606054
rect 3509 606051 3575 606054
rect 580165 604210 580231 604213
rect 583520 604210 584960 604300
rect 580165 604208 584960 604210
rect 580165 604152 580170 604208
rect 580226 604152 584960 604208
rect 580165 604150 584960 604152
rect 580165 604147 580231 604150
rect 583520 604060 584960 604150
rect 9397 596186 9463 596189
rect 9397 596184 12052 596186
rect 9397 596128 9402 596184
rect 9458 596128 12052 596184
rect 9397 596126 12052 596128
rect 9397 596123 9463 596126
rect 569309 595506 569375 595509
rect 566076 595504 569375 595506
rect 566076 595448 569314 595504
rect 569370 595448 569375 595504
rect 566076 595446 569375 595448
rect 569309 595443 569375 595446
rect -960 593058 480 593148
rect 2773 593058 2839 593061
rect -960 593056 2839 593058
rect -960 593000 2778 593056
rect 2834 593000 2839 593056
rect -960 592998 2839 593000
rect -960 592908 480 592998
rect 2773 592995 2839 592998
rect 579797 591018 579863 591021
rect 583520 591018 584960 591108
rect 579797 591016 584960 591018
rect 579797 590960 579802 591016
rect 579858 590960 584960 591016
rect 579797 590958 584960 590960
rect 579797 590955 579863 590958
rect 583520 590868 584960 590958
rect 9397 583946 9463 583949
rect 9397 583944 12052 583946
rect 9397 583888 9402 583944
rect 9458 583888 12052 583944
rect 9397 583886 12052 583888
rect 9397 583883 9463 583886
rect 569401 582994 569467 582997
rect 566076 582992 569467 582994
rect 566076 582936 569406 582992
rect 569462 582936 569467 582992
rect 566076 582934 569467 582936
rect 569401 582931 569467 582934
rect -960 580002 480 580092
rect 2957 580002 3023 580005
rect -960 580000 3023 580002
rect -960 579944 2962 580000
rect 3018 579944 3023 580000
rect -960 579942 3023 579944
rect -960 579852 480 579942
rect 2957 579939 3023 579942
rect 580165 577690 580231 577693
rect 583520 577690 584960 577780
rect 580165 577688 584960 577690
rect 580165 577632 580170 577688
rect 580226 577632 584960 577688
rect 580165 577630 584960 577632
rect 580165 577627 580231 577630
rect 583520 577540 584960 577630
rect 8845 571706 8911 571709
rect 8845 571704 12052 571706
rect 8845 571648 8850 571704
rect 8906 571648 12052 571704
rect 8845 571646 12052 571648
rect 8845 571643 8911 571646
rect 569217 570482 569283 570485
rect 566076 570480 569283 570482
rect 566076 570424 569222 570480
rect 569278 570424 569283 570480
rect 566076 570422 569283 570424
rect 569217 570419 569283 570422
rect -960 566946 480 567036
rect 3417 566946 3483 566949
rect -960 566944 3483 566946
rect -960 566888 3422 566944
rect 3478 566888 3483 566944
rect -960 566886 3483 566888
rect -960 566796 480 566886
rect 3417 566883 3483 566886
rect 579797 564362 579863 564365
rect 583520 564362 584960 564452
rect 579797 564360 584960 564362
rect 579797 564304 579802 564360
rect 579858 564304 584960 564360
rect 579797 564302 584960 564304
rect 579797 564299 579863 564302
rect 583520 564212 584960 564302
rect 9397 559466 9463 559469
rect 9397 559464 12052 559466
rect 9397 559408 9402 559464
rect 9458 559408 12052 559464
rect 9397 559406 12052 559408
rect 9397 559403 9463 559406
rect 569309 557970 569375 557973
rect 566076 557968 569375 557970
rect 566076 557912 569314 557968
rect 569370 557912 569375 557968
rect 566076 557910 569375 557912
rect 569309 557907 569375 557910
rect -960 553890 480 553980
rect 3509 553890 3575 553893
rect -960 553888 3575 553890
rect -960 553832 3514 553888
rect 3570 553832 3575 553888
rect -960 553830 3575 553832
rect -960 553740 480 553830
rect 3509 553827 3575 553830
rect 580165 551170 580231 551173
rect 583520 551170 584960 551260
rect 580165 551168 584960 551170
rect 580165 551112 580170 551168
rect 580226 551112 584960 551168
rect 580165 551110 584960 551112
rect 580165 551107 580231 551110
rect 583520 551020 584960 551110
rect 9397 547226 9463 547229
rect 9397 547224 12052 547226
rect 9397 547168 9402 547224
rect 9458 547168 12052 547224
rect 9397 547166 12052 547168
rect 9397 547163 9463 547166
rect 569217 545458 569283 545461
rect 566076 545456 569283 545458
rect 566076 545400 569222 545456
rect 569278 545400 569283 545456
rect 566076 545398 569283 545400
rect 569217 545395 569283 545398
rect -960 540834 480 540924
rect 3417 540834 3483 540837
rect -960 540832 3483 540834
rect -960 540776 3422 540832
rect 3478 540776 3483 540832
rect -960 540774 3483 540776
rect -960 540684 480 540774
rect 3417 540771 3483 540774
rect 580165 537842 580231 537845
rect 583520 537842 584960 537932
rect 580165 537840 584960 537842
rect 580165 537784 580170 537840
rect 580226 537784 584960 537840
rect 580165 537782 584960 537784
rect 580165 537779 580231 537782
rect 583520 537692 584960 537782
rect 9397 534986 9463 534989
rect 9397 534984 12052 534986
rect 9397 534928 9402 534984
rect 9458 534928 12052 534984
rect 9397 534926 12052 534928
rect 9397 534923 9463 534926
rect 569309 532946 569375 532949
rect 566076 532944 569375 532946
rect 566076 532888 569314 532944
rect 569370 532888 569375 532944
rect 566076 532886 569375 532888
rect 569309 532883 569375 532886
rect -960 527914 480 528004
rect 3417 527914 3483 527917
rect -960 527912 3483 527914
rect -960 527856 3422 527912
rect 3478 527856 3483 527912
rect -960 527854 3483 527856
rect -960 527764 480 527854
rect 3417 527851 3483 527854
rect 580165 524514 580231 524517
rect 583520 524514 584960 524604
rect 580165 524512 584960 524514
rect 580165 524456 580170 524512
rect 580226 524456 584960 524512
rect 580165 524454 584960 524456
rect 580165 524451 580231 524454
rect 583520 524364 584960 524454
rect 7649 522746 7715 522749
rect 7649 522744 12052 522746
rect 7649 522688 7654 522744
rect 7710 522688 12052 522744
rect 7649 522686 12052 522688
rect 7649 522683 7715 522686
rect 569217 520434 569283 520437
rect 566076 520432 569283 520434
rect 566076 520376 569222 520432
rect 569278 520376 569283 520432
rect 566076 520374 569283 520376
rect 569217 520371 569283 520374
rect -960 514858 480 514948
rect 3417 514858 3483 514861
rect -960 514856 3483 514858
rect -960 514800 3422 514856
rect 3478 514800 3483 514856
rect -960 514798 3483 514800
rect -960 514708 480 514798
rect 3417 514795 3483 514798
rect 580165 511322 580231 511325
rect 583520 511322 584960 511412
rect 580165 511320 584960 511322
rect 580165 511264 580170 511320
rect 580226 511264 584960 511320
rect 580165 511262 584960 511264
rect 580165 511259 580231 511262
rect 583520 511172 584960 511262
rect 7557 510506 7623 510509
rect 7557 510504 12052 510506
rect 7557 510448 7562 510504
rect 7618 510448 12052 510504
rect 7557 510446 12052 510448
rect 7557 510443 7623 510446
rect 569309 507922 569375 507925
rect 566076 507920 569375 507922
rect 566076 507864 569314 507920
rect 569370 507864 569375 507920
rect 566076 507862 569375 507864
rect 569309 507859 569375 507862
rect -960 501802 480 501892
rect 3049 501802 3115 501805
rect -960 501800 3115 501802
rect -960 501744 3054 501800
rect 3110 501744 3115 501800
rect -960 501742 3115 501744
rect -960 501652 480 501742
rect 3049 501739 3115 501742
rect 8937 498266 9003 498269
rect 8937 498264 12052 498266
rect 8937 498208 8942 498264
rect 8998 498208 12052 498264
rect 8937 498206 12052 498208
rect 8937 498203 9003 498206
rect 579889 497994 579955 497997
rect 583520 497994 584960 498084
rect 579889 497992 584960 497994
rect 579889 497936 579894 497992
rect 579950 497936 584960 497992
rect 579889 497934 584960 497936
rect 579889 497931 579955 497934
rect 583520 497844 584960 497934
rect 569217 495410 569283 495413
rect 566076 495408 569283 495410
rect 566076 495352 569222 495408
rect 569278 495352 569283 495408
rect 566076 495350 569283 495352
rect 569217 495347 569283 495350
rect -960 488746 480 488836
rect 3417 488746 3483 488749
rect -960 488744 3483 488746
rect -960 488688 3422 488744
rect 3478 488688 3483 488744
rect -960 488686 3483 488688
rect -960 488596 480 488686
rect 3417 488683 3483 488686
rect 9029 486026 9095 486029
rect 9029 486024 12052 486026
rect 9029 485968 9034 486024
rect 9090 485968 12052 486024
rect 9029 485966 12052 485968
rect 9029 485963 9095 485966
rect 580625 484666 580691 484669
rect 583520 484666 584960 484756
rect 580625 484664 584960 484666
rect 580625 484608 580630 484664
rect 580686 484608 584960 484664
rect 580625 484606 584960 484608
rect 580625 484603 580691 484606
rect 583520 484516 584960 484606
rect 569861 482898 569927 482901
rect 566076 482896 569927 482898
rect 566076 482840 569866 482896
rect 569922 482840 569927 482896
rect 566076 482838 569927 482840
rect 569861 482835 569927 482838
rect -960 475690 480 475780
rect 3417 475690 3483 475693
rect -960 475688 3483 475690
rect -960 475632 3422 475688
rect 3478 475632 3483 475688
rect -960 475630 3483 475632
rect -960 475540 480 475630
rect 3417 475627 3483 475630
rect 8937 473786 9003 473789
rect 8937 473784 12052 473786
rect 8937 473728 8942 473784
rect 8998 473728 12052 473784
rect 8937 473726 12052 473728
rect 8937 473723 9003 473726
rect 579981 471474 580047 471477
rect 583520 471474 584960 471564
rect 579981 471472 584960 471474
rect 579981 471416 579986 471472
rect 580042 471416 584960 471472
rect 579981 471414 584960 471416
rect 579981 471411 580047 471414
rect 583520 471324 584960 471414
rect 569861 470386 569927 470389
rect 566076 470384 569927 470386
rect 566076 470328 569866 470384
rect 569922 470328 569927 470384
rect 566076 470326 569927 470328
rect 569861 470323 569927 470326
rect -960 462634 480 462724
rect 3417 462634 3483 462637
rect -960 462632 3483 462634
rect -960 462576 3422 462632
rect 3478 462576 3483 462632
rect -960 462574 3483 462576
rect -960 462484 480 462574
rect 3417 462571 3483 462574
rect 9029 461546 9095 461549
rect 9029 461544 12052 461546
rect 9029 461488 9034 461544
rect 9090 461488 12052 461544
rect 9029 461486 12052 461488
rect 9029 461483 9095 461486
rect 580257 458146 580323 458149
rect 583520 458146 584960 458236
rect 580257 458144 584960 458146
rect 580257 458088 580262 458144
rect 580318 458088 584960 458144
rect 580257 458086 584960 458088
rect 580257 458083 580323 458086
rect 583520 457996 584960 458086
rect 569861 457874 569927 457877
rect 566076 457872 569927 457874
rect 566076 457816 569866 457872
rect 569922 457816 569927 457872
rect 566076 457814 569927 457816
rect 569861 457811 569927 457814
rect -960 449578 480 449668
rect 2773 449578 2839 449581
rect -960 449576 2839 449578
rect -960 449520 2778 449576
rect 2834 449520 2839 449576
rect -960 449518 2839 449520
rect -960 449428 480 449518
rect 2773 449515 2839 449518
rect 8937 449306 9003 449309
rect 8937 449304 12052 449306
rect 8937 449248 8942 449304
rect 8998 449248 12052 449304
rect 8937 449246 12052 449248
rect 8937 449243 9003 449246
rect 569125 445362 569191 445365
rect 566076 445360 569191 445362
rect 566076 445304 569130 445360
rect 569186 445304 569191 445360
rect 566076 445302 569191 445304
rect 569125 445299 569191 445302
rect 580349 444818 580415 444821
rect 583520 444818 584960 444908
rect 580349 444816 584960 444818
rect 580349 444760 580354 444816
rect 580410 444760 584960 444816
rect 580349 444758 584960 444760
rect 580349 444755 580415 444758
rect 583520 444668 584960 444758
rect 9397 437066 9463 437069
rect 9397 437064 12052 437066
rect 9397 437008 9402 437064
rect 9458 437008 12052 437064
rect 9397 437006 12052 437008
rect 9397 437003 9463 437006
rect -960 436658 480 436748
rect 2957 436658 3023 436661
rect -960 436656 3023 436658
rect -960 436600 2962 436656
rect 3018 436600 3023 436656
rect -960 436598 3023 436600
rect -960 436508 480 436598
rect 2957 436595 3023 436598
rect 569309 432850 569375 432853
rect 566076 432848 569375 432850
rect 566076 432792 569314 432848
rect 569370 432792 569375 432848
rect 566076 432790 569375 432792
rect 569309 432787 569375 432790
rect 580165 431626 580231 431629
rect 583520 431626 584960 431716
rect 580165 431624 584960 431626
rect 580165 431568 580170 431624
rect 580226 431568 584960 431624
rect 580165 431566 584960 431568
rect 580165 431563 580231 431566
rect 583520 431476 584960 431566
rect 9397 424826 9463 424829
rect 9397 424824 12052 424826
rect 9397 424768 9402 424824
rect 9458 424768 12052 424824
rect 9397 424766 12052 424768
rect 9397 424763 9463 424766
rect -960 423602 480 423692
rect 3417 423602 3483 423605
rect -960 423600 3483 423602
rect -960 423544 3422 423600
rect 3478 423544 3483 423600
rect -960 423542 3483 423544
rect -960 423452 480 423542
rect 3417 423539 3483 423542
rect 569217 420338 569283 420341
rect 566076 420336 569283 420338
rect 566076 420280 569222 420336
rect 569278 420280 569283 420336
rect 566076 420278 569283 420280
rect 569217 420275 569283 420278
rect 580165 418298 580231 418301
rect 583520 418298 584960 418388
rect 580165 418296 584960 418298
rect 580165 418240 580170 418296
rect 580226 418240 584960 418296
rect 580165 418238 584960 418240
rect 580165 418235 580231 418238
rect 583520 418148 584960 418238
rect 7557 412586 7623 412589
rect 7557 412584 12052 412586
rect 7557 412528 7562 412584
rect 7618 412528 12052 412584
rect 7557 412526 12052 412528
rect 7557 412523 7623 412526
rect -960 410546 480 410636
rect 3141 410546 3207 410549
rect -960 410544 3207 410546
rect -960 410488 3146 410544
rect 3202 410488 3207 410544
rect -960 410486 3207 410488
rect -960 410396 480 410486
rect 3141 410483 3207 410486
rect 569217 407826 569283 407829
rect 566076 407824 569283 407826
rect 566076 407768 569222 407824
rect 569278 407768 569283 407824
rect 566076 407766 569283 407768
rect 569217 407763 569283 407766
rect 580165 404970 580231 404973
rect 583520 404970 584960 405060
rect 580165 404968 584960 404970
rect 580165 404912 580170 404968
rect 580226 404912 584960 404968
rect 580165 404910 584960 404912
rect 580165 404907 580231 404910
rect 583520 404820 584960 404910
rect 7557 400346 7623 400349
rect 7557 400344 12052 400346
rect 7557 400288 7562 400344
rect 7618 400288 12052 400344
rect 7557 400286 12052 400288
rect 7557 400283 7623 400286
rect -960 397490 480 397580
rect 3417 397490 3483 397493
rect -960 397488 3483 397490
rect -960 397432 3422 397488
rect 3478 397432 3483 397488
rect -960 397430 3483 397432
rect -960 397340 480 397430
rect 3417 397427 3483 397430
rect 569125 395314 569191 395317
rect 566076 395312 569191 395314
rect 566076 395256 569130 395312
rect 569186 395256 569191 395312
rect 566076 395254 569191 395256
rect 569125 395251 569191 395254
rect 578877 391778 578943 391781
rect 583520 391778 584960 391868
rect 578877 391776 584960 391778
rect 578877 391720 578882 391776
rect 578938 391720 584960 391776
rect 578877 391718 584960 391720
rect 578877 391715 578943 391718
rect 583520 391628 584960 391718
rect 7557 388106 7623 388109
rect 7557 388104 12052 388106
rect 7557 388048 7562 388104
rect 7618 388048 12052 388104
rect 7557 388046 12052 388048
rect 7557 388043 7623 388046
rect -960 384434 480 384524
rect 3417 384434 3483 384437
rect -960 384432 3483 384434
rect -960 384376 3422 384432
rect 3478 384376 3483 384432
rect -960 384374 3483 384376
rect -960 384284 480 384374
rect 3417 384371 3483 384374
rect 569861 382802 569927 382805
rect 566076 382800 569927 382802
rect 566076 382744 569866 382800
rect 569922 382744 569927 382800
rect 566076 382742 569927 382744
rect 569861 382739 569927 382742
rect 578877 378450 578943 378453
rect 583520 378450 584960 378540
rect 578877 378448 584960 378450
rect 578877 378392 578882 378448
rect 578938 378392 584960 378448
rect 578877 378390 584960 378392
rect 578877 378387 578943 378390
rect 583520 378300 584960 378390
rect 7557 375866 7623 375869
rect 7557 375864 12052 375866
rect 7557 375808 7562 375864
rect 7618 375808 12052 375864
rect 7557 375806 12052 375808
rect 7557 375803 7623 375806
rect -960 371378 480 371468
rect 3417 371378 3483 371381
rect -960 371376 3483 371378
rect -960 371320 3422 371376
rect 3478 371320 3483 371376
rect -960 371318 3483 371320
rect -960 371228 480 371318
rect 3417 371315 3483 371318
rect 569585 370290 569651 370293
rect 566076 370288 569651 370290
rect 566076 370232 569590 370288
rect 569646 370232 569651 370288
rect 566076 370230 569651 370232
rect 569585 370227 569651 370230
rect 579613 365122 579679 365125
rect 583520 365122 584960 365212
rect 579613 365120 584960 365122
rect 579613 365064 579618 365120
rect 579674 365064 584960 365120
rect 579613 365062 584960 365064
rect 579613 365059 579679 365062
rect 583520 364972 584960 365062
rect 7557 363626 7623 363629
rect 7557 363624 12052 363626
rect 7557 363568 7562 363624
rect 7618 363568 12052 363624
rect 7557 363566 12052 363568
rect 7557 363563 7623 363566
rect -960 358458 480 358548
rect 2773 358458 2839 358461
rect -960 358456 2839 358458
rect -960 358400 2778 358456
rect 2834 358400 2839 358456
rect -960 358398 2839 358400
rect -960 358308 480 358398
rect 2773 358395 2839 358398
rect 569677 357778 569743 357781
rect 566076 357776 569743 357778
rect 566076 357720 569682 357776
rect 569738 357720 569743 357776
rect 566076 357718 569743 357720
rect 569677 357715 569743 357718
rect 579521 351930 579587 351933
rect 583520 351930 584960 352020
rect 579521 351928 584960 351930
rect 579521 351872 579526 351928
rect 579582 351872 584960 351928
rect 579521 351870 584960 351872
rect 579521 351867 579587 351870
rect 583520 351780 584960 351870
rect 8661 351386 8727 351389
rect 8661 351384 12052 351386
rect 8661 351328 8666 351384
rect 8722 351328 12052 351384
rect 8661 351326 12052 351328
rect 8661 351323 8727 351326
rect -960 345402 480 345492
rect 4061 345402 4127 345405
rect -960 345400 4127 345402
rect -960 345344 4066 345400
rect 4122 345344 4127 345400
rect -960 345342 4127 345344
rect -960 345252 480 345342
rect 4061 345339 4127 345342
rect 569677 345266 569743 345269
rect 566076 345264 569743 345266
rect 566076 345208 569682 345264
rect 569738 345208 569743 345264
rect 566076 345206 569743 345208
rect 569677 345203 569743 345206
rect 9397 339146 9463 339149
rect 9397 339144 12052 339146
rect 9397 339088 9402 339144
rect 9458 339088 12052 339144
rect 9397 339086 12052 339088
rect 9397 339083 9463 339086
rect 580165 338602 580231 338605
rect 583520 338602 584960 338692
rect 580165 338600 584960 338602
rect 580165 338544 580170 338600
rect 580226 338544 584960 338600
rect 580165 338542 584960 338544
rect 580165 338539 580231 338542
rect 583520 338452 584960 338542
rect 569217 332754 569283 332757
rect 566076 332752 569283 332754
rect 566076 332696 569222 332752
rect 569278 332696 569283 332752
rect 566076 332694 569283 332696
rect 569217 332691 569283 332694
rect -960 332346 480 332436
rect 3049 332346 3115 332349
rect -960 332344 3115 332346
rect -960 332288 3054 332344
rect 3110 332288 3115 332344
rect -960 332286 3115 332288
rect -960 332196 480 332286
rect 3049 332283 3115 332286
rect 9397 326906 9463 326909
rect 9397 326904 12052 326906
rect 9397 326848 9402 326904
rect 9458 326848 12052 326904
rect 9397 326846 12052 326848
rect 9397 326843 9463 326846
rect 580165 325274 580231 325277
rect 583520 325274 584960 325364
rect 580165 325272 584960 325274
rect 580165 325216 580170 325272
rect 580226 325216 584960 325272
rect 580165 325214 584960 325216
rect 580165 325211 580231 325214
rect 583520 325124 584960 325214
rect 568665 320242 568731 320245
rect 566076 320240 568731 320242
rect 566076 320184 568670 320240
rect 568726 320184 568731 320240
rect 566076 320182 568731 320184
rect 568665 320179 568731 320182
rect -960 319290 480 319380
rect 3417 319290 3483 319293
rect -960 319288 3483 319290
rect -960 319232 3422 319288
rect 3478 319232 3483 319288
rect -960 319230 3483 319232
rect -960 319140 480 319230
rect 3417 319227 3483 319230
rect 9397 314666 9463 314669
rect 9397 314664 12052 314666
rect 9397 314608 9402 314664
rect 9458 314608 12052 314664
rect 9397 314606 12052 314608
rect 9397 314603 9463 314606
rect 580165 312082 580231 312085
rect 583520 312082 584960 312172
rect 580165 312080 584960 312082
rect 580165 312024 580170 312080
rect 580226 312024 584960 312080
rect 580165 312022 584960 312024
rect 580165 312019 580231 312022
rect 583520 311932 584960 312022
rect 568941 307730 569007 307733
rect 566076 307728 569007 307730
rect 566076 307672 568946 307728
rect 569002 307672 569007 307728
rect 566076 307670 569007 307672
rect 568941 307667 569007 307670
rect -960 306234 480 306324
rect 3417 306234 3483 306237
rect -960 306232 3483 306234
rect -960 306176 3422 306232
rect 3478 306176 3483 306232
rect -960 306174 3483 306176
rect -960 306084 480 306174
rect 3417 306171 3483 306174
rect 9397 302426 9463 302429
rect 9397 302424 12052 302426
rect 9397 302368 9402 302424
rect 9458 302368 12052 302424
rect 9397 302366 12052 302368
rect 9397 302363 9463 302366
rect 580349 298754 580415 298757
rect 583520 298754 584960 298844
rect 580349 298752 584960 298754
rect 580349 298696 580354 298752
rect 580410 298696 584960 298752
rect 580349 298694 584960 298696
rect 580349 298691 580415 298694
rect 583520 298604 584960 298694
rect 569861 295218 569927 295221
rect 566076 295216 569927 295218
rect 566076 295160 569866 295216
rect 569922 295160 569927 295216
rect 566076 295158 569927 295160
rect 569861 295155 569927 295158
rect -960 293178 480 293268
rect 3417 293178 3483 293181
rect -960 293176 3483 293178
rect -960 293120 3422 293176
rect 3478 293120 3483 293176
rect -960 293118 3483 293120
rect -960 293028 480 293118
rect 3417 293115 3483 293118
rect 9397 290186 9463 290189
rect 9397 290184 12052 290186
rect 9397 290128 9402 290184
rect 9458 290128 12052 290184
rect 9397 290126 12052 290128
rect 9397 290123 9463 290126
rect 580165 285426 580231 285429
rect 583520 285426 584960 285516
rect 580165 285424 584960 285426
rect 580165 285368 580170 285424
rect 580226 285368 584960 285424
rect 580165 285366 584960 285368
rect 580165 285363 580231 285366
rect 583520 285276 584960 285366
rect 569861 282706 569927 282709
rect 566076 282704 569927 282706
rect 566076 282648 569866 282704
rect 569922 282648 569927 282704
rect 566076 282646 569927 282648
rect 569861 282643 569927 282646
rect -960 280122 480 280212
rect 3417 280122 3483 280125
rect -960 280120 3483 280122
rect -960 280064 3422 280120
rect 3478 280064 3483 280120
rect -960 280062 3483 280064
rect -960 279972 480 280062
rect 3417 280059 3483 280062
rect 9213 277946 9279 277949
rect 9213 277944 12052 277946
rect 9213 277888 9218 277944
rect 9274 277888 12052 277944
rect 9213 277886 12052 277888
rect 9213 277883 9279 277886
rect 579797 272234 579863 272237
rect 583520 272234 584960 272324
rect 579797 272232 584960 272234
rect 579797 272176 579802 272232
rect 579858 272176 584960 272232
rect 579797 272174 584960 272176
rect 579797 272171 579863 272174
rect 583520 272084 584960 272174
rect 569309 270194 569375 270197
rect 566076 270192 569375 270194
rect 566076 270136 569314 270192
rect 569370 270136 569375 270192
rect 566076 270134 569375 270136
rect 569309 270131 569375 270134
rect -960 267202 480 267292
rect 3049 267202 3115 267205
rect -960 267200 3115 267202
rect -960 267144 3054 267200
rect 3110 267144 3115 267200
rect -960 267142 3115 267144
rect -960 267052 480 267142
rect 3049 267139 3115 267142
rect 9397 265706 9463 265709
rect 9397 265704 12052 265706
rect 9397 265648 9402 265704
rect 9458 265648 12052 265704
rect 9397 265646 12052 265648
rect 9397 265643 9463 265646
rect 579705 258906 579771 258909
rect 583520 258906 584960 258996
rect 579705 258904 584960 258906
rect 579705 258848 579710 258904
rect 579766 258848 584960 258904
rect 579705 258846 584960 258848
rect 579705 258843 579771 258846
rect 583520 258756 584960 258846
rect 569125 257682 569191 257685
rect 566076 257680 569191 257682
rect 566076 257624 569130 257680
rect 569186 257624 569191 257680
rect 566076 257622 569191 257624
rect 569125 257619 569191 257622
rect -960 254146 480 254236
rect 3417 254146 3483 254149
rect -960 254144 3483 254146
rect -960 254088 3422 254144
rect 3478 254088 3483 254144
rect -960 254086 3483 254088
rect -960 253996 480 254086
rect 3417 254083 3483 254086
rect 9397 253466 9463 253469
rect 9397 253464 12052 253466
rect 9397 253408 9402 253464
rect 9458 253408 12052 253464
rect 9397 253406 12052 253408
rect 9397 253403 9463 253406
rect 580165 245578 580231 245581
rect 583520 245578 584960 245668
rect 580165 245576 584960 245578
rect 580165 245520 580170 245576
rect 580226 245520 584960 245576
rect 580165 245518 584960 245520
rect 580165 245515 580231 245518
rect 583520 245428 584960 245518
rect 568665 245170 568731 245173
rect 566076 245168 568731 245170
rect 566076 245112 568670 245168
rect 568726 245112 568731 245168
rect 566076 245110 568731 245112
rect 568665 245107 568731 245110
rect 9397 241226 9463 241229
rect 9397 241224 12052 241226
rect -960 241090 480 241180
rect 9397 241168 9402 241224
rect 9458 241168 12052 241224
rect 9397 241166 12052 241168
rect 9397 241163 9463 241166
rect 3417 241090 3483 241093
rect -960 241088 3483 241090
rect -960 241032 3422 241088
rect 3478 241032 3483 241088
rect -960 241030 3483 241032
rect -960 240940 480 241030
rect 3417 241027 3483 241030
rect 569861 232658 569927 232661
rect 566076 232656 569927 232658
rect 566076 232600 569866 232656
rect 569922 232600 569927 232656
rect 566076 232598 569927 232600
rect 569861 232595 569927 232598
rect 580165 232386 580231 232389
rect 583520 232386 584960 232476
rect 580165 232384 584960 232386
rect 580165 232328 580170 232384
rect 580226 232328 584960 232384
rect 580165 232326 584960 232328
rect 580165 232323 580231 232326
rect 583520 232236 584960 232326
rect 8845 228986 8911 228989
rect 8845 228984 12052 228986
rect 8845 228928 8850 228984
rect 8906 228928 12052 228984
rect 8845 228926 12052 228928
rect 8845 228923 8911 228926
rect -960 228034 480 228124
rect 3417 228034 3483 228037
rect -960 228032 3483 228034
rect -960 227976 3422 228032
rect 3478 227976 3483 228032
rect -960 227974 3483 227976
rect -960 227884 480 227974
rect 3417 227971 3483 227974
rect 569493 220146 569559 220149
rect 566076 220144 569559 220146
rect 566076 220088 569498 220144
rect 569554 220088 569559 220144
rect 566076 220086 569559 220088
rect 569493 220083 569559 220086
rect 580441 219058 580507 219061
rect 583520 219058 584960 219148
rect 580441 219056 584960 219058
rect 580441 219000 580446 219056
rect 580502 219000 584960 219056
rect 580441 218998 584960 219000
rect 580441 218995 580507 218998
rect 583520 218908 584960 218998
rect 8201 216746 8267 216749
rect 8201 216744 12052 216746
rect 8201 216688 8206 216744
rect 8262 216688 12052 216744
rect 8201 216686 12052 216688
rect 8201 216683 8267 216686
rect -960 214978 480 215068
rect 3417 214978 3483 214981
rect -960 214976 3483 214978
rect -960 214920 3422 214976
rect 3478 214920 3483 214976
rect -960 214918 3483 214920
rect -960 214828 480 214918
rect 3417 214915 3483 214918
rect 569861 207634 569927 207637
rect 566076 207632 569927 207634
rect 566076 207576 569866 207632
rect 569922 207576 569927 207632
rect 566076 207574 569927 207576
rect 569861 207571 569927 207574
rect 579521 205730 579587 205733
rect 583520 205730 584960 205820
rect 579521 205728 584960 205730
rect 579521 205672 579526 205728
rect 579582 205672 584960 205728
rect 579521 205670 584960 205672
rect 579521 205667 579587 205670
rect 583520 205580 584960 205670
rect 8201 204506 8267 204509
rect 8201 204504 12052 204506
rect 8201 204448 8206 204504
rect 8262 204448 12052 204504
rect 8201 204446 12052 204448
rect 8201 204443 8267 204446
rect -960 201922 480 202012
rect 3325 201922 3391 201925
rect -960 201920 3391 201922
rect -960 201864 3330 201920
rect 3386 201864 3391 201920
rect -960 201862 3391 201864
rect -960 201772 480 201862
rect 3325 201859 3391 201862
rect 569309 195122 569375 195125
rect 566076 195120 569375 195122
rect 566076 195064 569314 195120
rect 569370 195064 569375 195120
rect 566076 195062 569375 195064
rect 569309 195059 569375 195062
rect 579521 192538 579587 192541
rect 583520 192538 584960 192628
rect 579521 192536 584960 192538
rect 579521 192480 579526 192536
rect 579582 192480 584960 192536
rect 579521 192478 584960 192480
rect 579521 192475 579587 192478
rect 583520 192388 584960 192478
rect 8201 192266 8267 192269
rect 8201 192264 12052 192266
rect 8201 192208 8206 192264
rect 8262 192208 12052 192264
rect 8201 192206 12052 192208
rect 8201 192203 8267 192206
rect -960 188866 480 188956
rect 3417 188866 3483 188869
rect -960 188864 3483 188866
rect -960 188808 3422 188864
rect 3478 188808 3483 188864
rect -960 188806 3483 188808
rect -960 188716 480 188806
rect 3417 188803 3483 188806
rect 569401 182610 569467 182613
rect 566076 182608 569467 182610
rect 566076 182552 569406 182608
rect 569462 182552 569467 182608
rect 566076 182550 569467 182552
rect 569401 182547 569467 182550
rect 8201 180026 8267 180029
rect 8201 180024 12052 180026
rect 8201 179968 8206 180024
rect 8262 179968 12052 180024
rect 8201 179966 12052 179968
rect 8201 179963 8267 179966
rect 580257 179210 580323 179213
rect 583520 179210 584960 179300
rect 580257 179208 584960 179210
rect 580257 179152 580262 179208
rect 580318 179152 584960 179208
rect 580257 179150 584960 179152
rect 580257 179147 580323 179150
rect 583520 179060 584960 179150
rect -960 175946 480 176036
rect 3417 175946 3483 175949
rect -960 175944 3483 175946
rect -960 175888 3422 175944
rect 3478 175888 3483 175944
rect -960 175886 3483 175888
rect -960 175796 480 175886
rect 3417 175883 3483 175886
rect 569861 170098 569927 170101
rect 566076 170096 569927 170098
rect 566076 170040 569866 170096
rect 569922 170040 569927 170096
rect 566076 170038 569927 170040
rect 569861 170035 569927 170038
rect 8201 167786 8267 167789
rect 8201 167784 12052 167786
rect 8201 167728 8206 167784
rect 8262 167728 12052 167784
rect 8201 167726 12052 167728
rect 8201 167723 8267 167726
rect 579981 165882 580047 165885
rect 583520 165882 584960 165972
rect 579981 165880 584960 165882
rect 579981 165824 579986 165880
rect 580042 165824 584960 165880
rect 579981 165822 584960 165824
rect 579981 165819 580047 165822
rect 583520 165732 584960 165822
rect -960 162890 480 162980
rect 3509 162890 3575 162893
rect -960 162888 3575 162890
rect -960 162832 3514 162888
rect 3570 162832 3575 162888
rect -960 162830 3575 162832
rect -960 162740 480 162830
rect 3509 162827 3575 162830
rect 569861 157586 569927 157589
rect 566076 157584 569927 157586
rect 566076 157528 569866 157584
rect 569922 157528 569927 157584
rect 566076 157526 569927 157528
rect 569861 157523 569927 157526
rect 8937 155546 9003 155549
rect 8937 155544 12052 155546
rect 8937 155488 8942 155544
rect 8998 155488 12052 155544
rect 8937 155486 12052 155488
rect 8937 155483 9003 155486
rect 579521 152690 579587 152693
rect 583520 152690 584960 152780
rect 579521 152688 584960 152690
rect 579521 152632 579526 152688
rect 579582 152632 584960 152688
rect 579521 152630 584960 152632
rect 579521 152627 579587 152630
rect 583520 152540 584960 152630
rect -960 149834 480 149924
rect 3417 149834 3483 149837
rect -960 149832 3483 149834
rect -960 149776 3422 149832
rect 3478 149776 3483 149832
rect -960 149774 3483 149776
rect -960 149684 480 149774
rect 3417 149771 3483 149774
rect 569861 145074 569927 145077
rect 566076 145072 569927 145074
rect 566076 145016 569866 145072
rect 569922 145016 569927 145072
rect 566076 145014 569927 145016
rect 569861 145011 569927 145014
rect 8293 143306 8359 143309
rect 8293 143304 12052 143306
rect 8293 143248 8298 143304
rect 8354 143248 12052 143304
rect 8293 143246 12052 143248
rect 8293 143243 8359 143246
rect 578877 139362 578943 139365
rect 583520 139362 584960 139452
rect 578877 139360 584960 139362
rect 578877 139304 578882 139360
rect 578938 139304 584960 139360
rect 578877 139302 584960 139304
rect 578877 139299 578943 139302
rect 583520 139212 584960 139302
rect -960 136778 480 136868
rect 3233 136778 3299 136781
rect -960 136776 3299 136778
rect -960 136720 3238 136776
rect 3294 136720 3299 136776
rect -960 136718 3299 136720
rect -960 136628 480 136718
rect 3233 136715 3299 136718
rect 569861 132562 569927 132565
rect 566076 132560 569927 132562
rect 566076 132504 569866 132560
rect 569922 132504 569927 132560
rect 566076 132502 569927 132504
rect 569861 132499 569927 132502
rect 9029 131066 9095 131069
rect 9029 131064 12052 131066
rect 9029 131008 9034 131064
rect 9090 131008 12052 131064
rect 9029 131006 12052 131008
rect 9029 131003 9095 131006
rect 579613 126034 579679 126037
rect 583520 126034 584960 126124
rect 579613 126032 584960 126034
rect 579613 125976 579618 126032
rect 579674 125976 584960 126032
rect 579613 125974 584960 125976
rect 579613 125971 579679 125974
rect 583520 125884 584960 125974
rect -960 123722 480 123812
rect 4061 123722 4127 123725
rect -960 123720 4127 123722
rect -960 123664 4066 123720
rect 4122 123664 4127 123720
rect -960 123662 4127 123664
rect -960 123572 480 123662
rect 4061 123659 4127 123662
rect 568665 120050 568731 120053
rect 566076 120048 568731 120050
rect 566076 119992 568670 120048
rect 568726 119992 568731 120048
rect 566076 119990 568731 119992
rect 568665 119987 568731 119990
rect 9397 118826 9463 118829
rect 9397 118824 12052 118826
rect 9397 118768 9402 118824
rect 9458 118768 12052 118824
rect 9397 118766 12052 118768
rect 9397 118763 9463 118766
rect 578877 112842 578943 112845
rect 583520 112842 584960 112932
rect 578877 112840 584960 112842
rect 578877 112784 578882 112840
rect 578938 112784 584960 112840
rect 578877 112782 584960 112784
rect 578877 112779 578943 112782
rect 583520 112692 584960 112782
rect -960 110666 480 110756
rect 2773 110666 2839 110669
rect -960 110664 2839 110666
rect -960 110608 2778 110664
rect 2834 110608 2839 110664
rect -960 110606 2839 110608
rect -960 110516 480 110606
rect 2773 110603 2839 110606
rect 569677 107538 569743 107541
rect 566076 107536 569743 107538
rect 566076 107480 569682 107536
rect 569738 107480 569743 107536
rect 566076 107478 569743 107480
rect 569677 107475 569743 107478
rect 9397 106586 9463 106589
rect 9397 106584 12052 106586
rect 9397 106528 9402 106584
rect 9458 106528 12052 106584
rect 9397 106526 12052 106528
rect 9397 106523 9463 106526
rect 578877 99514 578943 99517
rect 583520 99514 584960 99604
rect 578877 99512 584960 99514
rect 578877 99456 578882 99512
rect 578938 99456 584960 99512
rect 578877 99454 584960 99456
rect 578877 99451 578943 99454
rect 583520 99364 584960 99454
rect -960 97610 480 97700
rect 2773 97610 2839 97613
rect -960 97608 2839 97610
rect -960 97552 2778 97608
rect 2834 97552 2839 97608
rect -960 97550 2839 97552
rect -960 97460 480 97550
rect 2773 97547 2839 97550
rect 569677 95026 569743 95029
rect 566076 95024 569743 95026
rect 566076 94968 569682 95024
rect 569738 94968 569743 95024
rect 566076 94966 569743 94968
rect 569677 94963 569743 94966
rect 9397 94346 9463 94349
rect 9397 94344 12052 94346
rect 9397 94288 9402 94344
rect 9458 94288 12052 94344
rect 9397 94286 12052 94288
rect 9397 94283 9463 94286
rect 580165 86186 580231 86189
rect 583520 86186 584960 86276
rect 580165 86184 584960 86186
rect 580165 86128 580170 86184
rect 580226 86128 584960 86184
rect 580165 86126 584960 86128
rect 580165 86123 580231 86126
rect 583520 86036 584960 86126
rect -960 84690 480 84780
rect 2773 84690 2839 84693
rect -960 84688 2839 84690
rect -960 84632 2778 84688
rect 2834 84632 2839 84688
rect -960 84630 2839 84632
rect -960 84540 480 84630
rect 2773 84627 2839 84630
rect 569677 82514 569743 82517
rect 566076 82512 569743 82514
rect 566076 82456 569682 82512
rect 569738 82456 569743 82512
rect 566076 82454 569743 82456
rect 569677 82451 569743 82454
rect 8937 82106 9003 82109
rect 8937 82104 12052 82106
rect 8937 82048 8942 82104
rect 8998 82048 12052 82104
rect 8937 82046 12052 82048
rect 8937 82043 9003 82046
rect 578877 72994 578943 72997
rect 583520 72994 584960 73084
rect 578877 72992 584960 72994
rect 578877 72936 578882 72992
rect 578938 72936 584960 72992
rect 578877 72934 584960 72936
rect 578877 72931 578943 72934
rect 583520 72844 584960 72934
rect -960 71634 480 71724
rect 3417 71634 3483 71637
rect -960 71632 3483 71634
rect -960 71576 3422 71632
rect 3478 71576 3483 71632
rect -960 71574 3483 71576
rect -960 71484 480 71574
rect 3417 71571 3483 71574
rect 569585 70002 569651 70005
rect 566076 70000 569651 70002
rect 566076 69944 569590 70000
rect 569646 69944 569651 70000
rect 566076 69942 569651 69944
rect 569585 69939 569651 69942
rect 8937 69866 9003 69869
rect 8937 69864 12052 69866
rect 8937 69808 8942 69864
rect 8998 69808 12052 69864
rect 8937 69806 12052 69808
rect 8937 69803 9003 69806
rect 578877 59666 578943 59669
rect 583520 59666 584960 59756
rect 578877 59664 584960 59666
rect 578877 59608 578882 59664
rect 578938 59608 584960 59664
rect 578877 59606 584960 59608
rect 578877 59603 578943 59606
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect 3141 58578 3207 58581
rect -960 58576 3207 58578
rect -960 58520 3146 58576
rect 3202 58520 3207 58576
rect -960 58518 3207 58520
rect -960 58428 480 58518
rect 3141 58515 3207 58518
rect 8845 57626 8911 57629
rect 8845 57624 12052 57626
rect 8845 57568 8850 57624
rect 8906 57568 12052 57624
rect 8845 57566 12052 57568
rect 8845 57563 8911 57566
rect 569125 57490 569191 57493
rect 566076 57488 569191 57490
rect 566076 57432 569130 57488
rect 569186 57432 569191 57488
rect 566076 57430 569191 57432
rect 569125 57427 569191 57430
rect 580165 46338 580231 46341
rect 583520 46338 584960 46428
rect 580165 46336 584960 46338
rect 580165 46280 580170 46336
rect 580226 46280 584960 46336
rect 580165 46278 584960 46280
rect 580165 46275 580231 46278
rect 583520 46188 584960 46278
rect -960 45522 480 45612
rect 2773 45522 2839 45525
rect -960 45520 2839 45522
rect -960 45464 2778 45520
rect 2834 45464 2839 45520
rect -960 45462 2839 45464
rect -960 45372 480 45462
rect 2773 45459 2839 45462
rect 9397 45386 9463 45389
rect 9397 45384 12052 45386
rect 9397 45328 9402 45384
rect 9458 45328 12052 45384
rect 9397 45326 12052 45328
rect 9397 45323 9463 45326
rect 569861 44978 569927 44981
rect 566076 44976 569927 44978
rect 566076 44920 569866 44976
rect 569922 44920 569927 44976
rect 566076 44918 569927 44920
rect 569861 44915 569927 44918
rect 9029 33146 9095 33149
rect 578877 33146 578943 33149
rect 583520 33146 584960 33236
rect 9029 33144 12052 33146
rect 9029 33088 9034 33144
rect 9090 33088 12052 33144
rect 9029 33086 12052 33088
rect 578877 33144 584960 33146
rect 578877 33088 578882 33144
rect 578938 33088 584960 33144
rect 578877 33086 584960 33088
rect 9029 33083 9095 33086
rect 578877 33083 578943 33086
rect 583520 32996 584960 33086
rect -960 32466 480 32556
rect 2773 32466 2839 32469
rect 569493 32466 569559 32469
rect -960 32464 2839 32466
rect -960 32408 2778 32464
rect 2834 32408 2839 32464
rect -960 32406 2839 32408
rect 566076 32464 569559 32466
rect 566076 32408 569498 32464
rect 569554 32408 569559 32464
rect 566076 32406 569559 32408
rect -960 32316 480 32406
rect 2773 32403 2839 32406
rect 569493 32403 569559 32406
rect 8937 20906 9003 20909
rect 8937 20904 12052 20906
rect 8937 20848 8942 20904
rect 8998 20848 12052 20904
rect 8937 20846 12052 20848
rect 8937 20843 9003 20846
rect 569861 19954 569927 19957
rect 566076 19952 569927 19954
rect 566076 19896 569866 19952
rect 569922 19896 569927 19952
rect 566076 19894 569927 19896
rect 569861 19891 569927 19894
rect 578969 19818 579035 19821
rect 583520 19818 584960 19908
rect 578969 19816 584960 19818
rect 578969 19760 578974 19816
rect 579030 19760 584960 19816
rect 578969 19758 584960 19760
rect 578969 19755 579035 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 2773 19410 2839 19413
rect -960 19408 2839 19410
rect -960 19352 2778 19408
rect 2834 19352 2839 19408
rect -960 19350 2839 19352
rect -960 19260 480 19350
rect 2773 19347 2839 19350
rect 578877 6626 578943 6629
rect 583520 6626 584960 6716
rect 578877 6624 584960 6626
rect -960 6490 480 6580
rect 578877 6568 578882 6624
rect 578938 6568 584960 6624
rect 578877 6566 584960 6568
rect 578877 6563 578943 6566
rect 3417 6490 3483 6493
rect -960 6488 3483 6490
rect -960 6432 3422 6488
rect 3478 6432 3483 6488
rect 583520 6476 584960 6566
rect -960 6430 3483 6432
rect -960 6340 480 6430
rect 3417 6427 3483 6430
rect 546493 4042 546559 4045
rect 568021 4042 568087 4045
rect 546493 4040 568087 4042
rect 546493 3984 546498 4040
rect 546554 3984 568026 4040
rect 568082 3984 568087 4040
rect 546493 3982 568087 3984
rect 546493 3979 546559 3982
rect 568021 3979 568087 3982
rect 536097 3906 536163 3909
rect 556337 3906 556403 3909
rect 536097 3904 556403 3906
rect 536097 3848 536102 3904
rect 536158 3848 556342 3904
rect 556398 3848 556403 3904
rect 536097 3846 556403 3848
rect 536097 3843 536163 3846
rect 556337 3843 556403 3846
rect 532785 3770 532851 3773
rect 553761 3770 553827 3773
rect 532785 3768 553827 3770
rect 532785 3712 532790 3768
rect 532846 3712 553766 3768
rect 553822 3712 553827 3768
rect 532785 3710 553827 3712
rect 532785 3707 532851 3710
rect 553761 3707 553827 3710
rect 559005 3770 559071 3773
rect 582189 3770 582255 3773
rect 559005 3768 582255 3770
rect 559005 3712 559010 3768
rect 559066 3712 582194 3768
rect 582250 3712 582255 3768
rect 559005 3710 582255 3712
rect 559005 3707 559071 3710
rect 582189 3707 582255 3710
rect 543641 3634 543707 3637
rect 564433 3634 564499 3637
rect 543641 3632 564499 3634
rect 543641 3576 543646 3632
rect 543702 3576 564438 3632
rect 564494 3576 564499 3632
rect 543641 3574 564499 3576
rect 543641 3571 543707 3574
rect 564433 3571 564499 3574
rect 549345 3498 549411 3501
rect 571517 3498 571583 3501
rect 549345 3496 571583 3498
rect 549345 3440 549350 3496
rect 549406 3440 571522 3496
rect 571578 3440 571583 3496
rect 549345 3438 571583 3440
rect 549345 3435 549411 3438
rect 571517 3435 571583 3438
rect 525977 3362 526043 3365
rect 546677 3362 546743 3365
rect 525977 3360 546743 3362
rect 525977 3304 525982 3360
rect 526038 3304 546682 3360
rect 546738 3304 546743 3360
rect 525977 3302 546743 3304
rect 525977 3299 526043 3302
rect 546677 3299 546743 3302
rect 548057 3362 548123 3365
rect 570321 3362 570387 3365
rect 548057 3360 570387 3362
rect 548057 3304 548062 3360
rect 548118 3304 570326 3360
rect 570382 3304 570387 3360
rect 548057 3302 570387 3304
rect 548057 3299 548123 3302
rect 570321 3299 570387 3302
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 677494 -8106 711002
rect -8726 677258 -8694 677494
rect -8458 677258 -8374 677494
rect -8138 677258 -8106 677494
rect -8726 677174 -8106 677258
rect -8726 676938 -8694 677174
rect -8458 676938 -8374 677174
rect -8138 676938 -8106 677174
rect -8726 641494 -8106 676938
rect -8726 641258 -8694 641494
rect -8458 641258 -8374 641494
rect -8138 641258 -8106 641494
rect -8726 641174 -8106 641258
rect -8726 640938 -8694 641174
rect -8458 640938 -8374 641174
rect -8138 640938 -8106 641174
rect -8726 605494 -8106 640938
rect -8726 605258 -8694 605494
rect -8458 605258 -8374 605494
rect -8138 605258 -8106 605494
rect -8726 605174 -8106 605258
rect -8726 604938 -8694 605174
rect -8458 604938 -8374 605174
rect -8138 604938 -8106 605174
rect -8726 569494 -8106 604938
rect -8726 569258 -8694 569494
rect -8458 569258 -8374 569494
rect -8138 569258 -8106 569494
rect -8726 569174 -8106 569258
rect -8726 568938 -8694 569174
rect -8458 568938 -8374 569174
rect -8138 568938 -8106 569174
rect -8726 533494 -8106 568938
rect -8726 533258 -8694 533494
rect -8458 533258 -8374 533494
rect -8138 533258 -8106 533494
rect -8726 533174 -8106 533258
rect -8726 532938 -8694 533174
rect -8458 532938 -8374 533174
rect -8138 532938 -8106 533174
rect -8726 497494 -8106 532938
rect -8726 497258 -8694 497494
rect -8458 497258 -8374 497494
rect -8138 497258 -8106 497494
rect -8726 497174 -8106 497258
rect -8726 496938 -8694 497174
rect -8458 496938 -8374 497174
rect -8138 496938 -8106 497174
rect -8726 461494 -8106 496938
rect -8726 461258 -8694 461494
rect -8458 461258 -8374 461494
rect -8138 461258 -8106 461494
rect -8726 461174 -8106 461258
rect -8726 460938 -8694 461174
rect -8458 460938 -8374 461174
rect -8138 460938 -8106 461174
rect -8726 425494 -8106 460938
rect -8726 425258 -8694 425494
rect -8458 425258 -8374 425494
rect -8138 425258 -8106 425494
rect -8726 425174 -8106 425258
rect -8726 424938 -8694 425174
rect -8458 424938 -8374 425174
rect -8138 424938 -8106 425174
rect -8726 389494 -8106 424938
rect -8726 389258 -8694 389494
rect -8458 389258 -8374 389494
rect -8138 389258 -8106 389494
rect -8726 389174 -8106 389258
rect -8726 388938 -8694 389174
rect -8458 388938 -8374 389174
rect -8138 388938 -8106 389174
rect -8726 353494 -8106 388938
rect -8726 353258 -8694 353494
rect -8458 353258 -8374 353494
rect -8138 353258 -8106 353494
rect -8726 353174 -8106 353258
rect -8726 352938 -8694 353174
rect -8458 352938 -8374 353174
rect -8138 352938 -8106 353174
rect -8726 317494 -8106 352938
rect -8726 317258 -8694 317494
rect -8458 317258 -8374 317494
rect -8138 317258 -8106 317494
rect -8726 317174 -8106 317258
rect -8726 316938 -8694 317174
rect -8458 316938 -8374 317174
rect -8138 316938 -8106 317174
rect -8726 281494 -8106 316938
rect -8726 281258 -8694 281494
rect -8458 281258 -8374 281494
rect -8138 281258 -8106 281494
rect -8726 281174 -8106 281258
rect -8726 280938 -8694 281174
rect -8458 280938 -8374 281174
rect -8138 280938 -8106 281174
rect -8726 245494 -8106 280938
rect -8726 245258 -8694 245494
rect -8458 245258 -8374 245494
rect -8138 245258 -8106 245494
rect -8726 245174 -8106 245258
rect -8726 244938 -8694 245174
rect -8458 244938 -8374 245174
rect -8138 244938 -8106 245174
rect -8726 209494 -8106 244938
rect -8726 209258 -8694 209494
rect -8458 209258 -8374 209494
rect -8138 209258 -8106 209494
rect -8726 209174 -8106 209258
rect -8726 208938 -8694 209174
rect -8458 208938 -8374 209174
rect -8138 208938 -8106 209174
rect -8726 173494 -8106 208938
rect -8726 173258 -8694 173494
rect -8458 173258 -8374 173494
rect -8138 173258 -8106 173494
rect -8726 173174 -8106 173258
rect -8726 172938 -8694 173174
rect -8458 172938 -8374 173174
rect -8138 172938 -8106 173174
rect -8726 137494 -8106 172938
rect -8726 137258 -8694 137494
rect -8458 137258 -8374 137494
rect -8138 137258 -8106 137494
rect -8726 137174 -8106 137258
rect -8726 136938 -8694 137174
rect -8458 136938 -8374 137174
rect -8138 136938 -8106 137174
rect -8726 101494 -8106 136938
rect -8726 101258 -8694 101494
rect -8458 101258 -8374 101494
rect -8138 101258 -8106 101494
rect -8726 101174 -8106 101258
rect -8726 100938 -8694 101174
rect -8458 100938 -8374 101174
rect -8138 100938 -8106 101174
rect -8726 65494 -8106 100938
rect -8726 65258 -8694 65494
rect -8458 65258 -8374 65494
rect -8138 65258 -8106 65494
rect -8726 65174 -8106 65258
rect -8726 64938 -8694 65174
rect -8458 64938 -8374 65174
rect -8138 64938 -8106 65174
rect -8726 29494 -8106 64938
rect -8726 29258 -8694 29494
rect -8458 29258 -8374 29494
rect -8138 29258 -8106 29494
rect -8726 29174 -8106 29258
rect -8726 28938 -8694 29174
rect -8458 28938 -8374 29174
rect -8138 28938 -8106 29174
rect -8726 -7066 -8106 28938
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 673774 -7146 710042
rect -7766 673538 -7734 673774
rect -7498 673538 -7414 673774
rect -7178 673538 -7146 673774
rect -7766 673454 -7146 673538
rect -7766 673218 -7734 673454
rect -7498 673218 -7414 673454
rect -7178 673218 -7146 673454
rect -7766 637774 -7146 673218
rect -7766 637538 -7734 637774
rect -7498 637538 -7414 637774
rect -7178 637538 -7146 637774
rect -7766 637454 -7146 637538
rect -7766 637218 -7734 637454
rect -7498 637218 -7414 637454
rect -7178 637218 -7146 637454
rect -7766 601774 -7146 637218
rect -7766 601538 -7734 601774
rect -7498 601538 -7414 601774
rect -7178 601538 -7146 601774
rect -7766 601454 -7146 601538
rect -7766 601218 -7734 601454
rect -7498 601218 -7414 601454
rect -7178 601218 -7146 601454
rect -7766 565774 -7146 601218
rect -7766 565538 -7734 565774
rect -7498 565538 -7414 565774
rect -7178 565538 -7146 565774
rect -7766 565454 -7146 565538
rect -7766 565218 -7734 565454
rect -7498 565218 -7414 565454
rect -7178 565218 -7146 565454
rect -7766 529774 -7146 565218
rect -7766 529538 -7734 529774
rect -7498 529538 -7414 529774
rect -7178 529538 -7146 529774
rect -7766 529454 -7146 529538
rect -7766 529218 -7734 529454
rect -7498 529218 -7414 529454
rect -7178 529218 -7146 529454
rect -7766 493774 -7146 529218
rect -7766 493538 -7734 493774
rect -7498 493538 -7414 493774
rect -7178 493538 -7146 493774
rect -7766 493454 -7146 493538
rect -7766 493218 -7734 493454
rect -7498 493218 -7414 493454
rect -7178 493218 -7146 493454
rect -7766 457774 -7146 493218
rect -7766 457538 -7734 457774
rect -7498 457538 -7414 457774
rect -7178 457538 -7146 457774
rect -7766 457454 -7146 457538
rect -7766 457218 -7734 457454
rect -7498 457218 -7414 457454
rect -7178 457218 -7146 457454
rect -7766 421774 -7146 457218
rect -7766 421538 -7734 421774
rect -7498 421538 -7414 421774
rect -7178 421538 -7146 421774
rect -7766 421454 -7146 421538
rect -7766 421218 -7734 421454
rect -7498 421218 -7414 421454
rect -7178 421218 -7146 421454
rect -7766 385774 -7146 421218
rect -7766 385538 -7734 385774
rect -7498 385538 -7414 385774
rect -7178 385538 -7146 385774
rect -7766 385454 -7146 385538
rect -7766 385218 -7734 385454
rect -7498 385218 -7414 385454
rect -7178 385218 -7146 385454
rect -7766 349774 -7146 385218
rect -7766 349538 -7734 349774
rect -7498 349538 -7414 349774
rect -7178 349538 -7146 349774
rect -7766 349454 -7146 349538
rect -7766 349218 -7734 349454
rect -7498 349218 -7414 349454
rect -7178 349218 -7146 349454
rect -7766 313774 -7146 349218
rect -7766 313538 -7734 313774
rect -7498 313538 -7414 313774
rect -7178 313538 -7146 313774
rect -7766 313454 -7146 313538
rect -7766 313218 -7734 313454
rect -7498 313218 -7414 313454
rect -7178 313218 -7146 313454
rect -7766 277774 -7146 313218
rect -7766 277538 -7734 277774
rect -7498 277538 -7414 277774
rect -7178 277538 -7146 277774
rect -7766 277454 -7146 277538
rect -7766 277218 -7734 277454
rect -7498 277218 -7414 277454
rect -7178 277218 -7146 277454
rect -7766 241774 -7146 277218
rect -7766 241538 -7734 241774
rect -7498 241538 -7414 241774
rect -7178 241538 -7146 241774
rect -7766 241454 -7146 241538
rect -7766 241218 -7734 241454
rect -7498 241218 -7414 241454
rect -7178 241218 -7146 241454
rect -7766 205774 -7146 241218
rect -7766 205538 -7734 205774
rect -7498 205538 -7414 205774
rect -7178 205538 -7146 205774
rect -7766 205454 -7146 205538
rect -7766 205218 -7734 205454
rect -7498 205218 -7414 205454
rect -7178 205218 -7146 205454
rect -7766 169774 -7146 205218
rect -7766 169538 -7734 169774
rect -7498 169538 -7414 169774
rect -7178 169538 -7146 169774
rect -7766 169454 -7146 169538
rect -7766 169218 -7734 169454
rect -7498 169218 -7414 169454
rect -7178 169218 -7146 169454
rect -7766 133774 -7146 169218
rect -7766 133538 -7734 133774
rect -7498 133538 -7414 133774
rect -7178 133538 -7146 133774
rect -7766 133454 -7146 133538
rect -7766 133218 -7734 133454
rect -7498 133218 -7414 133454
rect -7178 133218 -7146 133454
rect -7766 97774 -7146 133218
rect -7766 97538 -7734 97774
rect -7498 97538 -7414 97774
rect -7178 97538 -7146 97774
rect -7766 97454 -7146 97538
rect -7766 97218 -7734 97454
rect -7498 97218 -7414 97454
rect -7178 97218 -7146 97454
rect -7766 61774 -7146 97218
rect -7766 61538 -7734 61774
rect -7498 61538 -7414 61774
rect -7178 61538 -7146 61774
rect -7766 61454 -7146 61538
rect -7766 61218 -7734 61454
rect -7498 61218 -7414 61454
rect -7178 61218 -7146 61454
rect -7766 25774 -7146 61218
rect -7766 25538 -7734 25774
rect -7498 25538 -7414 25774
rect -7178 25538 -7146 25774
rect -7766 25454 -7146 25538
rect -7766 25218 -7734 25454
rect -7498 25218 -7414 25454
rect -7178 25218 -7146 25454
rect -7766 -6106 -7146 25218
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 670054 -6186 709082
rect -6806 669818 -6774 670054
rect -6538 669818 -6454 670054
rect -6218 669818 -6186 670054
rect -6806 669734 -6186 669818
rect -6806 669498 -6774 669734
rect -6538 669498 -6454 669734
rect -6218 669498 -6186 669734
rect -6806 634054 -6186 669498
rect -6806 633818 -6774 634054
rect -6538 633818 -6454 634054
rect -6218 633818 -6186 634054
rect -6806 633734 -6186 633818
rect -6806 633498 -6774 633734
rect -6538 633498 -6454 633734
rect -6218 633498 -6186 633734
rect -6806 598054 -6186 633498
rect -6806 597818 -6774 598054
rect -6538 597818 -6454 598054
rect -6218 597818 -6186 598054
rect -6806 597734 -6186 597818
rect -6806 597498 -6774 597734
rect -6538 597498 -6454 597734
rect -6218 597498 -6186 597734
rect -6806 562054 -6186 597498
rect -6806 561818 -6774 562054
rect -6538 561818 -6454 562054
rect -6218 561818 -6186 562054
rect -6806 561734 -6186 561818
rect -6806 561498 -6774 561734
rect -6538 561498 -6454 561734
rect -6218 561498 -6186 561734
rect -6806 526054 -6186 561498
rect -6806 525818 -6774 526054
rect -6538 525818 -6454 526054
rect -6218 525818 -6186 526054
rect -6806 525734 -6186 525818
rect -6806 525498 -6774 525734
rect -6538 525498 -6454 525734
rect -6218 525498 -6186 525734
rect -6806 490054 -6186 525498
rect -6806 489818 -6774 490054
rect -6538 489818 -6454 490054
rect -6218 489818 -6186 490054
rect -6806 489734 -6186 489818
rect -6806 489498 -6774 489734
rect -6538 489498 -6454 489734
rect -6218 489498 -6186 489734
rect -6806 454054 -6186 489498
rect -6806 453818 -6774 454054
rect -6538 453818 -6454 454054
rect -6218 453818 -6186 454054
rect -6806 453734 -6186 453818
rect -6806 453498 -6774 453734
rect -6538 453498 -6454 453734
rect -6218 453498 -6186 453734
rect -6806 418054 -6186 453498
rect -6806 417818 -6774 418054
rect -6538 417818 -6454 418054
rect -6218 417818 -6186 418054
rect -6806 417734 -6186 417818
rect -6806 417498 -6774 417734
rect -6538 417498 -6454 417734
rect -6218 417498 -6186 417734
rect -6806 382054 -6186 417498
rect -6806 381818 -6774 382054
rect -6538 381818 -6454 382054
rect -6218 381818 -6186 382054
rect -6806 381734 -6186 381818
rect -6806 381498 -6774 381734
rect -6538 381498 -6454 381734
rect -6218 381498 -6186 381734
rect -6806 346054 -6186 381498
rect -6806 345818 -6774 346054
rect -6538 345818 -6454 346054
rect -6218 345818 -6186 346054
rect -6806 345734 -6186 345818
rect -6806 345498 -6774 345734
rect -6538 345498 -6454 345734
rect -6218 345498 -6186 345734
rect -6806 310054 -6186 345498
rect -6806 309818 -6774 310054
rect -6538 309818 -6454 310054
rect -6218 309818 -6186 310054
rect -6806 309734 -6186 309818
rect -6806 309498 -6774 309734
rect -6538 309498 -6454 309734
rect -6218 309498 -6186 309734
rect -6806 274054 -6186 309498
rect -6806 273818 -6774 274054
rect -6538 273818 -6454 274054
rect -6218 273818 -6186 274054
rect -6806 273734 -6186 273818
rect -6806 273498 -6774 273734
rect -6538 273498 -6454 273734
rect -6218 273498 -6186 273734
rect -6806 238054 -6186 273498
rect -6806 237818 -6774 238054
rect -6538 237818 -6454 238054
rect -6218 237818 -6186 238054
rect -6806 237734 -6186 237818
rect -6806 237498 -6774 237734
rect -6538 237498 -6454 237734
rect -6218 237498 -6186 237734
rect -6806 202054 -6186 237498
rect -6806 201818 -6774 202054
rect -6538 201818 -6454 202054
rect -6218 201818 -6186 202054
rect -6806 201734 -6186 201818
rect -6806 201498 -6774 201734
rect -6538 201498 -6454 201734
rect -6218 201498 -6186 201734
rect -6806 166054 -6186 201498
rect -6806 165818 -6774 166054
rect -6538 165818 -6454 166054
rect -6218 165818 -6186 166054
rect -6806 165734 -6186 165818
rect -6806 165498 -6774 165734
rect -6538 165498 -6454 165734
rect -6218 165498 -6186 165734
rect -6806 130054 -6186 165498
rect -6806 129818 -6774 130054
rect -6538 129818 -6454 130054
rect -6218 129818 -6186 130054
rect -6806 129734 -6186 129818
rect -6806 129498 -6774 129734
rect -6538 129498 -6454 129734
rect -6218 129498 -6186 129734
rect -6806 94054 -6186 129498
rect -6806 93818 -6774 94054
rect -6538 93818 -6454 94054
rect -6218 93818 -6186 94054
rect -6806 93734 -6186 93818
rect -6806 93498 -6774 93734
rect -6538 93498 -6454 93734
rect -6218 93498 -6186 93734
rect -6806 58054 -6186 93498
rect -6806 57818 -6774 58054
rect -6538 57818 -6454 58054
rect -6218 57818 -6186 58054
rect -6806 57734 -6186 57818
rect -6806 57498 -6774 57734
rect -6538 57498 -6454 57734
rect -6218 57498 -6186 57734
rect -6806 22054 -6186 57498
rect -6806 21818 -6774 22054
rect -6538 21818 -6454 22054
rect -6218 21818 -6186 22054
rect -6806 21734 -6186 21818
rect -6806 21498 -6774 21734
rect -6538 21498 -6454 21734
rect -6218 21498 -6186 21734
rect -6806 -5146 -6186 21498
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 666334 -5226 708122
rect -5846 666098 -5814 666334
rect -5578 666098 -5494 666334
rect -5258 666098 -5226 666334
rect -5846 666014 -5226 666098
rect -5846 665778 -5814 666014
rect -5578 665778 -5494 666014
rect -5258 665778 -5226 666014
rect -5846 630334 -5226 665778
rect -5846 630098 -5814 630334
rect -5578 630098 -5494 630334
rect -5258 630098 -5226 630334
rect -5846 630014 -5226 630098
rect -5846 629778 -5814 630014
rect -5578 629778 -5494 630014
rect -5258 629778 -5226 630014
rect -5846 594334 -5226 629778
rect -5846 594098 -5814 594334
rect -5578 594098 -5494 594334
rect -5258 594098 -5226 594334
rect -5846 594014 -5226 594098
rect -5846 593778 -5814 594014
rect -5578 593778 -5494 594014
rect -5258 593778 -5226 594014
rect -5846 558334 -5226 593778
rect -5846 558098 -5814 558334
rect -5578 558098 -5494 558334
rect -5258 558098 -5226 558334
rect -5846 558014 -5226 558098
rect -5846 557778 -5814 558014
rect -5578 557778 -5494 558014
rect -5258 557778 -5226 558014
rect -5846 522334 -5226 557778
rect -5846 522098 -5814 522334
rect -5578 522098 -5494 522334
rect -5258 522098 -5226 522334
rect -5846 522014 -5226 522098
rect -5846 521778 -5814 522014
rect -5578 521778 -5494 522014
rect -5258 521778 -5226 522014
rect -5846 486334 -5226 521778
rect -5846 486098 -5814 486334
rect -5578 486098 -5494 486334
rect -5258 486098 -5226 486334
rect -5846 486014 -5226 486098
rect -5846 485778 -5814 486014
rect -5578 485778 -5494 486014
rect -5258 485778 -5226 486014
rect -5846 450334 -5226 485778
rect -5846 450098 -5814 450334
rect -5578 450098 -5494 450334
rect -5258 450098 -5226 450334
rect -5846 450014 -5226 450098
rect -5846 449778 -5814 450014
rect -5578 449778 -5494 450014
rect -5258 449778 -5226 450014
rect -5846 414334 -5226 449778
rect -5846 414098 -5814 414334
rect -5578 414098 -5494 414334
rect -5258 414098 -5226 414334
rect -5846 414014 -5226 414098
rect -5846 413778 -5814 414014
rect -5578 413778 -5494 414014
rect -5258 413778 -5226 414014
rect -5846 378334 -5226 413778
rect -5846 378098 -5814 378334
rect -5578 378098 -5494 378334
rect -5258 378098 -5226 378334
rect -5846 378014 -5226 378098
rect -5846 377778 -5814 378014
rect -5578 377778 -5494 378014
rect -5258 377778 -5226 378014
rect -5846 342334 -5226 377778
rect -5846 342098 -5814 342334
rect -5578 342098 -5494 342334
rect -5258 342098 -5226 342334
rect -5846 342014 -5226 342098
rect -5846 341778 -5814 342014
rect -5578 341778 -5494 342014
rect -5258 341778 -5226 342014
rect -5846 306334 -5226 341778
rect -5846 306098 -5814 306334
rect -5578 306098 -5494 306334
rect -5258 306098 -5226 306334
rect -5846 306014 -5226 306098
rect -5846 305778 -5814 306014
rect -5578 305778 -5494 306014
rect -5258 305778 -5226 306014
rect -5846 270334 -5226 305778
rect -5846 270098 -5814 270334
rect -5578 270098 -5494 270334
rect -5258 270098 -5226 270334
rect -5846 270014 -5226 270098
rect -5846 269778 -5814 270014
rect -5578 269778 -5494 270014
rect -5258 269778 -5226 270014
rect -5846 234334 -5226 269778
rect -5846 234098 -5814 234334
rect -5578 234098 -5494 234334
rect -5258 234098 -5226 234334
rect -5846 234014 -5226 234098
rect -5846 233778 -5814 234014
rect -5578 233778 -5494 234014
rect -5258 233778 -5226 234014
rect -5846 198334 -5226 233778
rect -5846 198098 -5814 198334
rect -5578 198098 -5494 198334
rect -5258 198098 -5226 198334
rect -5846 198014 -5226 198098
rect -5846 197778 -5814 198014
rect -5578 197778 -5494 198014
rect -5258 197778 -5226 198014
rect -5846 162334 -5226 197778
rect -5846 162098 -5814 162334
rect -5578 162098 -5494 162334
rect -5258 162098 -5226 162334
rect -5846 162014 -5226 162098
rect -5846 161778 -5814 162014
rect -5578 161778 -5494 162014
rect -5258 161778 -5226 162014
rect -5846 126334 -5226 161778
rect -5846 126098 -5814 126334
rect -5578 126098 -5494 126334
rect -5258 126098 -5226 126334
rect -5846 126014 -5226 126098
rect -5846 125778 -5814 126014
rect -5578 125778 -5494 126014
rect -5258 125778 -5226 126014
rect -5846 90334 -5226 125778
rect -5846 90098 -5814 90334
rect -5578 90098 -5494 90334
rect -5258 90098 -5226 90334
rect -5846 90014 -5226 90098
rect -5846 89778 -5814 90014
rect -5578 89778 -5494 90014
rect -5258 89778 -5226 90014
rect -5846 54334 -5226 89778
rect -5846 54098 -5814 54334
rect -5578 54098 -5494 54334
rect -5258 54098 -5226 54334
rect -5846 54014 -5226 54098
rect -5846 53778 -5814 54014
rect -5578 53778 -5494 54014
rect -5258 53778 -5226 54014
rect -5846 18334 -5226 53778
rect -5846 18098 -5814 18334
rect -5578 18098 -5494 18334
rect -5258 18098 -5226 18334
rect -5846 18014 -5226 18098
rect -5846 17778 -5814 18014
rect -5578 17778 -5494 18014
rect -5258 17778 -5226 18014
rect -5846 -4186 -5226 17778
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 698614 -4266 707162
rect -4886 698378 -4854 698614
rect -4618 698378 -4534 698614
rect -4298 698378 -4266 698614
rect -4886 698294 -4266 698378
rect -4886 698058 -4854 698294
rect -4618 698058 -4534 698294
rect -4298 698058 -4266 698294
rect -4886 662614 -4266 698058
rect -4886 662378 -4854 662614
rect -4618 662378 -4534 662614
rect -4298 662378 -4266 662614
rect -4886 662294 -4266 662378
rect -4886 662058 -4854 662294
rect -4618 662058 -4534 662294
rect -4298 662058 -4266 662294
rect -4886 626614 -4266 662058
rect -4886 626378 -4854 626614
rect -4618 626378 -4534 626614
rect -4298 626378 -4266 626614
rect -4886 626294 -4266 626378
rect -4886 626058 -4854 626294
rect -4618 626058 -4534 626294
rect -4298 626058 -4266 626294
rect -4886 590614 -4266 626058
rect -4886 590378 -4854 590614
rect -4618 590378 -4534 590614
rect -4298 590378 -4266 590614
rect -4886 590294 -4266 590378
rect -4886 590058 -4854 590294
rect -4618 590058 -4534 590294
rect -4298 590058 -4266 590294
rect -4886 554614 -4266 590058
rect -4886 554378 -4854 554614
rect -4618 554378 -4534 554614
rect -4298 554378 -4266 554614
rect -4886 554294 -4266 554378
rect -4886 554058 -4854 554294
rect -4618 554058 -4534 554294
rect -4298 554058 -4266 554294
rect -4886 518614 -4266 554058
rect -4886 518378 -4854 518614
rect -4618 518378 -4534 518614
rect -4298 518378 -4266 518614
rect -4886 518294 -4266 518378
rect -4886 518058 -4854 518294
rect -4618 518058 -4534 518294
rect -4298 518058 -4266 518294
rect -4886 482614 -4266 518058
rect -4886 482378 -4854 482614
rect -4618 482378 -4534 482614
rect -4298 482378 -4266 482614
rect -4886 482294 -4266 482378
rect -4886 482058 -4854 482294
rect -4618 482058 -4534 482294
rect -4298 482058 -4266 482294
rect -4886 446614 -4266 482058
rect -4886 446378 -4854 446614
rect -4618 446378 -4534 446614
rect -4298 446378 -4266 446614
rect -4886 446294 -4266 446378
rect -4886 446058 -4854 446294
rect -4618 446058 -4534 446294
rect -4298 446058 -4266 446294
rect -4886 410614 -4266 446058
rect -4886 410378 -4854 410614
rect -4618 410378 -4534 410614
rect -4298 410378 -4266 410614
rect -4886 410294 -4266 410378
rect -4886 410058 -4854 410294
rect -4618 410058 -4534 410294
rect -4298 410058 -4266 410294
rect -4886 374614 -4266 410058
rect -4886 374378 -4854 374614
rect -4618 374378 -4534 374614
rect -4298 374378 -4266 374614
rect -4886 374294 -4266 374378
rect -4886 374058 -4854 374294
rect -4618 374058 -4534 374294
rect -4298 374058 -4266 374294
rect -4886 338614 -4266 374058
rect -4886 338378 -4854 338614
rect -4618 338378 -4534 338614
rect -4298 338378 -4266 338614
rect -4886 338294 -4266 338378
rect -4886 338058 -4854 338294
rect -4618 338058 -4534 338294
rect -4298 338058 -4266 338294
rect -4886 302614 -4266 338058
rect -4886 302378 -4854 302614
rect -4618 302378 -4534 302614
rect -4298 302378 -4266 302614
rect -4886 302294 -4266 302378
rect -4886 302058 -4854 302294
rect -4618 302058 -4534 302294
rect -4298 302058 -4266 302294
rect -4886 266614 -4266 302058
rect -4886 266378 -4854 266614
rect -4618 266378 -4534 266614
rect -4298 266378 -4266 266614
rect -4886 266294 -4266 266378
rect -4886 266058 -4854 266294
rect -4618 266058 -4534 266294
rect -4298 266058 -4266 266294
rect -4886 230614 -4266 266058
rect -4886 230378 -4854 230614
rect -4618 230378 -4534 230614
rect -4298 230378 -4266 230614
rect -4886 230294 -4266 230378
rect -4886 230058 -4854 230294
rect -4618 230058 -4534 230294
rect -4298 230058 -4266 230294
rect -4886 194614 -4266 230058
rect -4886 194378 -4854 194614
rect -4618 194378 -4534 194614
rect -4298 194378 -4266 194614
rect -4886 194294 -4266 194378
rect -4886 194058 -4854 194294
rect -4618 194058 -4534 194294
rect -4298 194058 -4266 194294
rect -4886 158614 -4266 194058
rect -4886 158378 -4854 158614
rect -4618 158378 -4534 158614
rect -4298 158378 -4266 158614
rect -4886 158294 -4266 158378
rect -4886 158058 -4854 158294
rect -4618 158058 -4534 158294
rect -4298 158058 -4266 158294
rect -4886 122614 -4266 158058
rect -4886 122378 -4854 122614
rect -4618 122378 -4534 122614
rect -4298 122378 -4266 122614
rect -4886 122294 -4266 122378
rect -4886 122058 -4854 122294
rect -4618 122058 -4534 122294
rect -4298 122058 -4266 122294
rect -4886 86614 -4266 122058
rect -4886 86378 -4854 86614
rect -4618 86378 -4534 86614
rect -4298 86378 -4266 86614
rect -4886 86294 -4266 86378
rect -4886 86058 -4854 86294
rect -4618 86058 -4534 86294
rect -4298 86058 -4266 86294
rect -4886 50614 -4266 86058
rect -4886 50378 -4854 50614
rect -4618 50378 -4534 50614
rect -4298 50378 -4266 50614
rect -4886 50294 -4266 50378
rect -4886 50058 -4854 50294
rect -4618 50058 -4534 50294
rect -4298 50058 -4266 50294
rect -4886 14614 -4266 50058
rect -4886 14378 -4854 14614
rect -4618 14378 -4534 14614
rect -4298 14378 -4266 14614
rect -4886 14294 -4266 14378
rect -4886 14058 -4854 14294
rect -4618 14058 -4534 14294
rect -4298 14058 -4266 14294
rect -4886 -3226 -4266 14058
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 694894 -3306 706202
rect -3926 694658 -3894 694894
rect -3658 694658 -3574 694894
rect -3338 694658 -3306 694894
rect -3926 694574 -3306 694658
rect -3926 694338 -3894 694574
rect -3658 694338 -3574 694574
rect -3338 694338 -3306 694574
rect -3926 658894 -3306 694338
rect -3926 658658 -3894 658894
rect -3658 658658 -3574 658894
rect -3338 658658 -3306 658894
rect -3926 658574 -3306 658658
rect -3926 658338 -3894 658574
rect -3658 658338 -3574 658574
rect -3338 658338 -3306 658574
rect -3926 622894 -3306 658338
rect -3926 622658 -3894 622894
rect -3658 622658 -3574 622894
rect -3338 622658 -3306 622894
rect -3926 622574 -3306 622658
rect -3926 622338 -3894 622574
rect -3658 622338 -3574 622574
rect -3338 622338 -3306 622574
rect -3926 586894 -3306 622338
rect -3926 586658 -3894 586894
rect -3658 586658 -3574 586894
rect -3338 586658 -3306 586894
rect -3926 586574 -3306 586658
rect -3926 586338 -3894 586574
rect -3658 586338 -3574 586574
rect -3338 586338 -3306 586574
rect -3926 550894 -3306 586338
rect -3926 550658 -3894 550894
rect -3658 550658 -3574 550894
rect -3338 550658 -3306 550894
rect -3926 550574 -3306 550658
rect -3926 550338 -3894 550574
rect -3658 550338 -3574 550574
rect -3338 550338 -3306 550574
rect -3926 514894 -3306 550338
rect -3926 514658 -3894 514894
rect -3658 514658 -3574 514894
rect -3338 514658 -3306 514894
rect -3926 514574 -3306 514658
rect -3926 514338 -3894 514574
rect -3658 514338 -3574 514574
rect -3338 514338 -3306 514574
rect -3926 478894 -3306 514338
rect -3926 478658 -3894 478894
rect -3658 478658 -3574 478894
rect -3338 478658 -3306 478894
rect -3926 478574 -3306 478658
rect -3926 478338 -3894 478574
rect -3658 478338 -3574 478574
rect -3338 478338 -3306 478574
rect -3926 442894 -3306 478338
rect -3926 442658 -3894 442894
rect -3658 442658 -3574 442894
rect -3338 442658 -3306 442894
rect -3926 442574 -3306 442658
rect -3926 442338 -3894 442574
rect -3658 442338 -3574 442574
rect -3338 442338 -3306 442574
rect -3926 406894 -3306 442338
rect -3926 406658 -3894 406894
rect -3658 406658 -3574 406894
rect -3338 406658 -3306 406894
rect -3926 406574 -3306 406658
rect -3926 406338 -3894 406574
rect -3658 406338 -3574 406574
rect -3338 406338 -3306 406574
rect -3926 370894 -3306 406338
rect -3926 370658 -3894 370894
rect -3658 370658 -3574 370894
rect -3338 370658 -3306 370894
rect -3926 370574 -3306 370658
rect -3926 370338 -3894 370574
rect -3658 370338 -3574 370574
rect -3338 370338 -3306 370574
rect -3926 334894 -3306 370338
rect -3926 334658 -3894 334894
rect -3658 334658 -3574 334894
rect -3338 334658 -3306 334894
rect -3926 334574 -3306 334658
rect -3926 334338 -3894 334574
rect -3658 334338 -3574 334574
rect -3338 334338 -3306 334574
rect -3926 298894 -3306 334338
rect -3926 298658 -3894 298894
rect -3658 298658 -3574 298894
rect -3338 298658 -3306 298894
rect -3926 298574 -3306 298658
rect -3926 298338 -3894 298574
rect -3658 298338 -3574 298574
rect -3338 298338 -3306 298574
rect -3926 262894 -3306 298338
rect -3926 262658 -3894 262894
rect -3658 262658 -3574 262894
rect -3338 262658 -3306 262894
rect -3926 262574 -3306 262658
rect -3926 262338 -3894 262574
rect -3658 262338 -3574 262574
rect -3338 262338 -3306 262574
rect -3926 226894 -3306 262338
rect -3926 226658 -3894 226894
rect -3658 226658 -3574 226894
rect -3338 226658 -3306 226894
rect -3926 226574 -3306 226658
rect -3926 226338 -3894 226574
rect -3658 226338 -3574 226574
rect -3338 226338 -3306 226574
rect -3926 190894 -3306 226338
rect -3926 190658 -3894 190894
rect -3658 190658 -3574 190894
rect -3338 190658 -3306 190894
rect -3926 190574 -3306 190658
rect -3926 190338 -3894 190574
rect -3658 190338 -3574 190574
rect -3338 190338 -3306 190574
rect -3926 154894 -3306 190338
rect -3926 154658 -3894 154894
rect -3658 154658 -3574 154894
rect -3338 154658 -3306 154894
rect -3926 154574 -3306 154658
rect -3926 154338 -3894 154574
rect -3658 154338 -3574 154574
rect -3338 154338 -3306 154574
rect -3926 118894 -3306 154338
rect -3926 118658 -3894 118894
rect -3658 118658 -3574 118894
rect -3338 118658 -3306 118894
rect -3926 118574 -3306 118658
rect -3926 118338 -3894 118574
rect -3658 118338 -3574 118574
rect -3338 118338 -3306 118574
rect -3926 82894 -3306 118338
rect -3926 82658 -3894 82894
rect -3658 82658 -3574 82894
rect -3338 82658 -3306 82894
rect -3926 82574 -3306 82658
rect -3926 82338 -3894 82574
rect -3658 82338 -3574 82574
rect -3338 82338 -3306 82574
rect -3926 46894 -3306 82338
rect -3926 46658 -3894 46894
rect -3658 46658 -3574 46894
rect -3338 46658 -3306 46894
rect -3926 46574 -3306 46658
rect -3926 46338 -3894 46574
rect -3658 46338 -3574 46574
rect -3338 46338 -3306 46574
rect -3926 10894 -3306 46338
rect -3926 10658 -3894 10894
rect -3658 10658 -3574 10894
rect -3338 10658 -3306 10894
rect -3926 10574 -3306 10658
rect -3926 10338 -3894 10574
rect -3658 10338 -3574 10574
rect -3338 10338 -3306 10574
rect -3926 -2266 -3306 10338
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 691174 -2346 705242
rect -2966 690938 -2934 691174
rect -2698 690938 -2614 691174
rect -2378 690938 -2346 691174
rect -2966 690854 -2346 690938
rect -2966 690618 -2934 690854
rect -2698 690618 -2614 690854
rect -2378 690618 -2346 690854
rect -2966 655174 -2346 690618
rect -2966 654938 -2934 655174
rect -2698 654938 -2614 655174
rect -2378 654938 -2346 655174
rect -2966 654854 -2346 654938
rect -2966 654618 -2934 654854
rect -2698 654618 -2614 654854
rect -2378 654618 -2346 654854
rect -2966 619174 -2346 654618
rect -2966 618938 -2934 619174
rect -2698 618938 -2614 619174
rect -2378 618938 -2346 619174
rect -2966 618854 -2346 618938
rect -2966 618618 -2934 618854
rect -2698 618618 -2614 618854
rect -2378 618618 -2346 618854
rect -2966 583174 -2346 618618
rect -2966 582938 -2934 583174
rect -2698 582938 -2614 583174
rect -2378 582938 -2346 583174
rect -2966 582854 -2346 582938
rect -2966 582618 -2934 582854
rect -2698 582618 -2614 582854
rect -2378 582618 -2346 582854
rect -2966 547174 -2346 582618
rect -2966 546938 -2934 547174
rect -2698 546938 -2614 547174
rect -2378 546938 -2346 547174
rect -2966 546854 -2346 546938
rect -2966 546618 -2934 546854
rect -2698 546618 -2614 546854
rect -2378 546618 -2346 546854
rect -2966 511174 -2346 546618
rect -2966 510938 -2934 511174
rect -2698 510938 -2614 511174
rect -2378 510938 -2346 511174
rect -2966 510854 -2346 510938
rect -2966 510618 -2934 510854
rect -2698 510618 -2614 510854
rect -2378 510618 -2346 510854
rect -2966 475174 -2346 510618
rect -2966 474938 -2934 475174
rect -2698 474938 -2614 475174
rect -2378 474938 -2346 475174
rect -2966 474854 -2346 474938
rect -2966 474618 -2934 474854
rect -2698 474618 -2614 474854
rect -2378 474618 -2346 474854
rect -2966 439174 -2346 474618
rect -2966 438938 -2934 439174
rect -2698 438938 -2614 439174
rect -2378 438938 -2346 439174
rect -2966 438854 -2346 438938
rect -2966 438618 -2934 438854
rect -2698 438618 -2614 438854
rect -2378 438618 -2346 438854
rect -2966 403174 -2346 438618
rect -2966 402938 -2934 403174
rect -2698 402938 -2614 403174
rect -2378 402938 -2346 403174
rect -2966 402854 -2346 402938
rect -2966 402618 -2934 402854
rect -2698 402618 -2614 402854
rect -2378 402618 -2346 402854
rect -2966 367174 -2346 402618
rect -2966 366938 -2934 367174
rect -2698 366938 -2614 367174
rect -2378 366938 -2346 367174
rect -2966 366854 -2346 366938
rect -2966 366618 -2934 366854
rect -2698 366618 -2614 366854
rect -2378 366618 -2346 366854
rect -2966 331174 -2346 366618
rect -2966 330938 -2934 331174
rect -2698 330938 -2614 331174
rect -2378 330938 -2346 331174
rect -2966 330854 -2346 330938
rect -2966 330618 -2934 330854
rect -2698 330618 -2614 330854
rect -2378 330618 -2346 330854
rect -2966 295174 -2346 330618
rect -2966 294938 -2934 295174
rect -2698 294938 -2614 295174
rect -2378 294938 -2346 295174
rect -2966 294854 -2346 294938
rect -2966 294618 -2934 294854
rect -2698 294618 -2614 294854
rect -2378 294618 -2346 294854
rect -2966 259174 -2346 294618
rect -2966 258938 -2934 259174
rect -2698 258938 -2614 259174
rect -2378 258938 -2346 259174
rect -2966 258854 -2346 258938
rect -2966 258618 -2934 258854
rect -2698 258618 -2614 258854
rect -2378 258618 -2346 258854
rect -2966 223174 -2346 258618
rect -2966 222938 -2934 223174
rect -2698 222938 -2614 223174
rect -2378 222938 -2346 223174
rect -2966 222854 -2346 222938
rect -2966 222618 -2934 222854
rect -2698 222618 -2614 222854
rect -2378 222618 -2346 222854
rect -2966 187174 -2346 222618
rect -2966 186938 -2934 187174
rect -2698 186938 -2614 187174
rect -2378 186938 -2346 187174
rect -2966 186854 -2346 186938
rect -2966 186618 -2934 186854
rect -2698 186618 -2614 186854
rect -2378 186618 -2346 186854
rect -2966 151174 -2346 186618
rect -2966 150938 -2934 151174
rect -2698 150938 -2614 151174
rect -2378 150938 -2346 151174
rect -2966 150854 -2346 150938
rect -2966 150618 -2934 150854
rect -2698 150618 -2614 150854
rect -2378 150618 -2346 150854
rect -2966 115174 -2346 150618
rect -2966 114938 -2934 115174
rect -2698 114938 -2614 115174
rect -2378 114938 -2346 115174
rect -2966 114854 -2346 114938
rect -2966 114618 -2934 114854
rect -2698 114618 -2614 114854
rect -2378 114618 -2346 114854
rect -2966 79174 -2346 114618
rect -2966 78938 -2934 79174
rect -2698 78938 -2614 79174
rect -2378 78938 -2346 79174
rect -2966 78854 -2346 78938
rect -2966 78618 -2934 78854
rect -2698 78618 -2614 78854
rect -2378 78618 -2346 78854
rect -2966 43174 -2346 78618
rect -2966 42938 -2934 43174
rect -2698 42938 -2614 43174
rect -2378 42938 -2346 43174
rect -2966 42854 -2346 42938
rect -2966 42618 -2934 42854
rect -2698 42618 -2614 42854
rect -2378 42618 -2346 42854
rect -2966 7174 -2346 42618
rect -2966 6938 -2934 7174
rect -2698 6938 -2614 7174
rect -2378 6938 -2346 7174
rect -2966 6854 -2346 6938
rect -2966 6618 -2934 6854
rect -2698 6618 -2614 6854
rect -2378 6618 -2346 6854
rect -2966 -1306 -2346 6618
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 711590
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 1794 -7654 2414 -902
rect 5514 705798 6134 711590
rect 5514 705562 5546 705798
rect 5782 705562 5866 705798
rect 6102 705562 6134 705798
rect 5514 705478 6134 705562
rect 5514 705242 5546 705478
rect 5782 705242 5866 705478
rect 6102 705242 6134 705478
rect 5514 691174 6134 705242
rect 5514 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 6134 691174
rect 5514 690854 6134 690938
rect 5514 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 6134 690854
rect 5514 655174 6134 690618
rect 5514 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 6134 655174
rect 5514 654854 6134 654938
rect 5514 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 6134 654854
rect 5514 619174 6134 654618
rect 5514 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 6134 619174
rect 5514 618854 6134 618938
rect 5514 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 6134 618854
rect 5514 583174 6134 618618
rect 5514 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 6134 583174
rect 5514 582854 6134 582938
rect 5514 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 6134 582854
rect 5514 547174 6134 582618
rect 5514 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 6134 547174
rect 5514 546854 6134 546938
rect 5514 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 6134 546854
rect 5514 511174 6134 546618
rect 5514 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 6134 511174
rect 5514 510854 6134 510938
rect 5514 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 6134 510854
rect 5514 475174 6134 510618
rect 5514 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 6134 475174
rect 5514 474854 6134 474938
rect 5514 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 6134 474854
rect 5514 439174 6134 474618
rect 5514 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 6134 439174
rect 5514 438854 6134 438938
rect 5514 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 6134 438854
rect 5514 403174 6134 438618
rect 5514 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 6134 403174
rect 5514 402854 6134 402938
rect 5514 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 6134 402854
rect 5514 367174 6134 402618
rect 5514 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 6134 367174
rect 5514 366854 6134 366938
rect 5514 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 6134 366854
rect 5514 331174 6134 366618
rect 5514 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 6134 331174
rect 5514 330854 6134 330938
rect 5514 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 6134 330854
rect 5514 295174 6134 330618
rect 5514 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 6134 295174
rect 5514 294854 6134 294938
rect 5514 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 6134 294854
rect 5514 259174 6134 294618
rect 5514 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 6134 259174
rect 5514 258854 6134 258938
rect 5514 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 6134 258854
rect 5514 223174 6134 258618
rect 5514 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 6134 223174
rect 5514 222854 6134 222938
rect 5514 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 6134 222854
rect 5514 187174 6134 222618
rect 5514 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 6134 187174
rect 5514 186854 6134 186938
rect 5514 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 6134 186854
rect 5514 151174 6134 186618
rect 5514 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 6134 151174
rect 5514 150854 6134 150938
rect 5514 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 6134 150854
rect 5514 115174 6134 150618
rect 5514 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 6134 115174
rect 5514 114854 6134 114938
rect 5514 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 6134 114854
rect 5514 79174 6134 114618
rect 5514 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 6134 79174
rect 5514 78854 6134 78938
rect 5514 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 6134 78854
rect 5514 43174 6134 78618
rect 5514 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 6134 43174
rect 5514 42854 6134 42938
rect 5514 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 6134 42854
rect 5514 7174 6134 42618
rect 5514 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 6134 7174
rect 5514 6854 6134 6938
rect 5514 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 6134 6854
rect 5514 -1306 6134 6618
rect 5514 -1542 5546 -1306
rect 5782 -1542 5866 -1306
rect 6102 -1542 6134 -1306
rect 5514 -1626 6134 -1542
rect 5514 -1862 5546 -1626
rect 5782 -1862 5866 -1626
rect 6102 -1862 6134 -1626
rect 5514 -7654 6134 -1862
rect 9234 706758 9854 711590
rect 9234 706522 9266 706758
rect 9502 706522 9586 706758
rect 9822 706522 9854 706758
rect 9234 706438 9854 706522
rect 9234 706202 9266 706438
rect 9502 706202 9586 706438
rect 9822 706202 9854 706438
rect 9234 694894 9854 706202
rect 9234 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 9854 694894
rect 9234 694574 9854 694658
rect 9234 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 9854 694574
rect 9234 658894 9854 694338
rect 12954 707718 13574 711590
rect 12954 707482 12986 707718
rect 13222 707482 13306 707718
rect 13542 707482 13574 707718
rect 12954 707398 13574 707482
rect 12954 707162 12986 707398
rect 13222 707162 13306 707398
rect 13542 707162 13574 707398
rect 12954 698614 13574 707162
rect 12954 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 13574 698614
rect 12954 698294 13574 698378
rect 12954 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 13574 698294
rect 12954 677977 13574 698058
rect 37794 704838 38414 711590
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 677977 38414 686898
rect 41514 705798 42134 711590
rect 41514 705562 41546 705798
rect 41782 705562 41866 705798
rect 42102 705562 42134 705798
rect 41514 705478 42134 705562
rect 41514 705242 41546 705478
rect 41782 705242 41866 705478
rect 42102 705242 42134 705478
rect 41514 691174 42134 705242
rect 41514 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 42134 691174
rect 41514 690854 42134 690938
rect 41514 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 42134 690854
rect 41514 677977 42134 690618
rect 45234 706758 45854 711590
rect 45234 706522 45266 706758
rect 45502 706522 45586 706758
rect 45822 706522 45854 706758
rect 45234 706438 45854 706522
rect 45234 706202 45266 706438
rect 45502 706202 45586 706438
rect 45822 706202 45854 706438
rect 45234 694894 45854 706202
rect 45234 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 45854 694894
rect 45234 694574 45854 694658
rect 45234 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 45854 694574
rect 45234 677977 45854 694338
rect 48954 707718 49574 711590
rect 48954 707482 48986 707718
rect 49222 707482 49306 707718
rect 49542 707482 49574 707718
rect 48954 707398 49574 707482
rect 48954 707162 48986 707398
rect 49222 707162 49306 707398
rect 49542 707162 49574 707398
rect 48954 698614 49574 707162
rect 48954 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 49574 698614
rect 48954 698294 49574 698378
rect 48954 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 49574 698294
rect 48954 677977 49574 698058
rect 73794 704838 74414 711590
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 677977 74414 686898
rect 77514 705798 78134 711590
rect 77514 705562 77546 705798
rect 77782 705562 77866 705798
rect 78102 705562 78134 705798
rect 77514 705478 78134 705562
rect 77514 705242 77546 705478
rect 77782 705242 77866 705478
rect 78102 705242 78134 705478
rect 77514 691174 78134 705242
rect 77514 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 78134 691174
rect 77514 690854 78134 690938
rect 77514 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 78134 690854
rect 77514 678332 78134 690618
rect 81234 706758 81854 711590
rect 81234 706522 81266 706758
rect 81502 706522 81586 706758
rect 81822 706522 81854 706758
rect 81234 706438 81854 706522
rect 81234 706202 81266 706438
rect 81502 706202 81586 706438
rect 81822 706202 81854 706438
rect 81234 694894 81854 706202
rect 81234 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 81854 694894
rect 81234 694574 81854 694658
rect 81234 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 81854 694574
rect 81234 677977 81854 694338
rect 84954 707718 85574 711590
rect 84954 707482 84986 707718
rect 85222 707482 85306 707718
rect 85542 707482 85574 707718
rect 84954 707398 85574 707482
rect 84954 707162 84986 707398
rect 85222 707162 85306 707398
rect 85542 707162 85574 707398
rect 84954 698614 85574 707162
rect 84954 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 85574 698614
rect 84954 698294 85574 698378
rect 84954 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 85574 698294
rect 84954 677977 85574 698058
rect 109794 704838 110414 711590
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 677977 110414 686898
rect 113514 705798 114134 711590
rect 113514 705562 113546 705798
rect 113782 705562 113866 705798
rect 114102 705562 114134 705798
rect 113514 705478 114134 705562
rect 113514 705242 113546 705478
rect 113782 705242 113866 705478
rect 114102 705242 114134 705478
rect 113514 691174 114134 705242
rect 113514 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 114134 691174
rect 113514 690854 114134 690938
rect 113514 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 114134 690854
rect 113514 677977 114134 690618
rect 117234 706758 117854 711590
rect 117234 706522 117266 706758
rect 117502 706522 117586 706758
rect 117822 706522 117854 706758
rect 117234 706438 117854 706522
rect 117234 706202 117266 706438
rect 117502 706202 117586 706438
rect 117822 706202 117854 706438
rect 117234 694894 117854 706202
rect 117234 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 117854 694894
rect 117234 694574 117854 694658
rect 117234 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 117854 694574
rect 117234 677977 117854 694338
rect 120954 707718 121574 711590
rect 120954 707482 120986 707718
rect 121222 707482 121306 707718
rect 121542 707482 121574 707718
rect 120954 707398 121574 707482
rect 120954 707162 120986 707398
rect 121222 707162 121306 707398
rect 121542 707162 121574 707398
rect 120954 698614 121574 707162
rect 120954 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 121574 698614
rect 120954 698294 121574 698378
rect 120954 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 121574 698294
rect 120954 677977 121574 698058
rect 145794 704838 146414 711590
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 677977 146414 686898
rect 149514 705798 150134 711590
rect 149514 705562 149546 705798
rect 149782 705562 149866 705798
rect 150102 705562 150134 705798
rect 149514 705478 150134 705562
rect 149514 705242 149546 705478
rect 149782 705242 149866 705478
rect 150102 705242 150134 705478
rect 149514 691174 150134 705242
rect 149514 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 150134 691174
rect 149514 690854 150134 690938
rect 149514 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 150134 690854
rect 149514 677977 150134 690618
rect 153234 706758 153854 711590
rect 153234 706522 153266 706758
rect 153502 706522 153586 706758
rect 153822 706522 153854 706758
rect 153234 706438 153854 706522
rect 153234 706202 153266 706438
rect 153502 706202 153586 706438
rect 153822 706202 153854 706438
rect 153234 694894 153854 706202
rect 153234 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 153854 694894
rect 153234 694574 153854 694658
rect 153234 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 153854 694574
rect 153234 677977 153854 694338
rect 156954 707718 157574 711590
rect 156954 707482 156986 707718
rect 157222 707482 157306 707718
rect 157542 707482 157574 707718
rect 156954 707398 157574 707482
rect 156954 707162 156986 707398
rect 157222 707162 157306 707398
rect 157542 707162 157574 707398
rect 156954 698614 157574 707162
rect 156954 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 157574 698614
rect 156954 698294 157574 698378
rect 156954 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 157574 698294
rect 156954 677977 157574 698058
rect 181794 704838 182414 711590
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 677977 182414 686898
rect 185514 705798 186134 711590
rect 185514 705562 185546 705798
rect 185782 705562 185866 705798
rect 186102 705562 186134 705798
rect 185514 705478 186134 705562
rect 185514 705242 185546 705478
rect 185782 705242 185866 705478
rect 186102 705242 186134 705478
rect 185514 691174 186134 705242
rect 185514 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 186134 691174
rect 185514 690854 186134 690938
rect 185514 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 186134 690854
rect 185514 678332 186134 690618
rect 189234 706758 189854 711590
rect 189234 706522 189266 706758
rect 189502 706522 189586 706758
rect 189822 706522 189854 706758
rect 189234 706438 189854 706522
rect 189234 706202 189266 706438
rect 189502 706202 189586 706438
rect 189822 706202 189854 706438
rect 189234 694894 189854 706202
rect 189234 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 189854 694894
rect 189234 694574 189854 694658
rect 189234 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 189854 694574
rect 189234 677977 189854 694338
rect 192954 707718 193574 711590
rect 192954 707482 192986 707718
rect 193222 707482 193306 707718
rect 193542 707482 193574 707718
rect 192954 707398 193574 707482
rect 192954 707162 192986 707398
rect 193222 707162 193306 707398
rect 193542 707162 193574 707398
rect 192954 698614 193574 707162
rect 192954 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 193574 698614
rect 192954 698294 193574 698378
rect 192954 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 193574 698294
rect 192954 677977 193574 698058
rect 217794 704838 218414 711590
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 677977 218414 686898
rect 221514 705798 222134 711590
rect 221514 705562 221546 705798
rect 221782 705562 221866 705798
rect 222102 705562 222134 705798
rect 221514 705478 222134 705562
rect 221514 705242 221546 705478
rect 221782 705242 221866 705478
rect 222102 705242 222134 705478
rect 221514 691174 222134 705242
rect 221514 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 222134 691174
rect 221514 690854 222134 690938
rect 221514 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 222134 690854
rect 221514 677977 222134 690618
rect 225234 706758 225854 711590
rect 225234 706522 225266 706758
rect 225502 706522 225586 706758
rect 225822 706522 225854 706758
rect 225234 706438 225854 706522
rect 225234 706202 225266 706438
rect 225502 706202 225586 706438
rect 225822 706202 225854 706438
rect 225234 694894 225854 706202
rect 225234 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 225854 694894
rect 225234 694574 225854 694658
rect 225234 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 225854 694574
rect 225234 677977 225854 694338
rect 228954 707718 229574 711590
rect 228954 707482 228986 707718
rect 229222 707482 229306 707718
rect 229542 707482 229574 707718
rect 228954 707398 229574 707482
rect 228954 707162 228986 707398
rect 229222 707162 229306 707398
rect 229542 707162 229574 707398
rect 228954 698614 229574 707162
rect 228954 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 229574 698614
rect 228954 698294 229574 698378
rect 228954 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 229574 698294
rect 228954 677977 229574 698058
rect 253794 704838 254414 711590
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 677977 254414 686898
rect 257514 705798 258134 711590
rect 257514 705562 257546 705798
rect 257782 705562 257866 705798
rect 258102 705562 258134 705798
rect 257514 705478 258134 705562
rect 257514 705242 257546 705478
rect 257782 705242 257866 705478
rect 258102 705242 258134 705478
rect 257514 691174 258134 705242
rect 257514 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 258134 691174
rect 257514 690854 258134 690938
rect 257514 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 258134 690854
rect 257514 677977 258134 690618
rect 261234 706758 261854 711590
rect 261234 706522 261266 706758
rect 261502 706522 261586 706758
rect 261822 706522 261854 706758
rect 261234 706438 261854 706522
rect 261234 706202 261266 706438
rect 261502 706202 261586 706438
rect 261822 706202 261854 706438
rect 261234 694894 261854 706202
rect 261234 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 261854 694894
rect 261234 694574 261854 694658
rect 261234 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 261854 694574
rect 261234 677977 261854 694338
rect 264954 707718 265574 711590
rect 264954 707482 264986 707718
rect 265222 707482 265306 707718
rect 265542 707482 265574 707718
rect 264954 707398 265574 707482
rect 264954 707162 264986 707398
rect 265222 707162 265306 707398
rect 265542 707162 265574 707398
rect 264954 698614 265574 707162
rect 264954 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 265574 698614
rect 264954 698294 265574 698378
rect 264954 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 265574 698294
rect 264954 677977 265574 698058
rect 289794 704838 290414 711590
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 677977 290414 686898
rect 293514 705798 294134 711590
rect 293514 705562 293546 705798
rect 293782 705562 293866 705798
rect 294102 705562 294134 705798
rect 293514 705478 294134 705562
rect 293514 705242 293546 705478
rect 293782 705242 293866 705478
rect 294102 705242 294134 705478
rect 293514 691174 294134 705242
rect 293514 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 294134 691174
rect 293514 690854 294134 690938
rect 293514 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 294134 690854
rect 293514 677977 294134 690618
rect 297234 706758 297854 711590
rect 297234 706522 297266 706758
rect 297502 706522 297586 706758
rect 297822 706522 297854 706758
rect 297234 706438 297854 706522
rect 297234 706202 297266 706438
rect 297502 706202 297586 706438
rect 297822 706202 297854 706438
rect 297234 694894 297854 706202
rect 297234 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 297854 694894
rect 297234 694574 297854 694658
rect 297234 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 297854 694574
rect 297234 677977 297854 694338
rect 300954 707718 301574 711590
rect 300954 707482 300986 707718
rect 301222 707482 301306 707718
rect 301542 707482 301574 707718
rect 300954 707398 301574 707482
rect 300954 707162 300986 707398
rect 301222 707162 301306 707398
rect 301542 707162 301574 707398
rect 300954 698614 301574 707162
rect 300954 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 301574 698614
rect 300954 698294 301574 698378
rect 300954 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 301574 698294
rect 300954 677977 301574 698058
rect 325794 704838 326414 711590
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 677977 326414 686898
rect 329514 705798 330134 711590
rect 329514 705562 329546 705798
rect 329782 705562 329866 705798
rect 330102 705562 330134 705798
rect 329514 705478 330134 705562
rect 329514 705242 329546 705478
rect 329782 705242 329866 705478
rect 330102 705242 330134 705478
rect 329514 691174 330134 705242
rect 329514 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 330134 691174
rect 329514 690854 330134 690938
rect 329514 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 330134 690854
rect 329514 677977 330134 690618
rect 333234 706758 333854 711590
rect 333234 706522 333266 706758
rect 333502 706522 333586 706758
rect 333822 706522 333854 706758
rect 333234 706438 333854 706522
rect 333234 706202 333266 706438
rect 333502 706202 333586 706438
rect 333822 706202 333854 706438
rect 333234 694894 333854 706202
rect 333234 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 333854 694894
rect 333234 694574 333854 694658
rect 333234 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 333854 694574
rect 333234 677977 333854 694338
rect 336954 707718 337574 711590
rect 336954 707482 336986 707718
rect 337222 707482 337306 707718
rect 337542 707482 337574 707718
rect 336954 707398 337574 707482
rect 336954 707162 336986 707398
rect 337222 707162 337306 707398
rect 337542 707162 337574 707398
rect 336954 698614 337574 707162
rect 336954 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 337574 698614
rect 336954 698294 337574 698378
rect 336954 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 337574 698294
rect 336954 677977 337574 698058
rect 361794 704838 362414 711590
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 677977 362414 686898
rect 365514 705798 366134 711590
rect 365514 705562 365546 705798
rect 365782 705562 365866 705798
rect 366102 705562 366134 705798
rect 365514 705478 366134 705562
rect 365514 705242 365546 705478
rect 365782 705242 365866 705478
rect 366102 705242 366134 705478
rect 365514 691174 366134 705242
rect 365514 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 366134 691174
rect 365514 690854 366134 690938
rect 365514 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 366134 690854
rect 365514 677977 366134 690618
rect 369234 706758 369854 711590
rect 369234 706522 369266 706758
rect 369502 706522 369586 706758
rect 369822 706522 369854 706758
rect 369234 706438 369854 706522
rect 369234 706202 369266 706438
rect 369502 706202 369586 706438
rect 369822 706202 369854 706438
rect 369234 694894 369854 706202
rect 369234 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 369854 694894
rect 369234 694574 369854 694658
rect 369234 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 369854 694574
rect 369234 678332 369854 694338
rect 372954 707718 373574 711590
rect 372954 707482 372986 707718
rect 373222 707482 373306 707718
rect 373542 707482 373574 707718
rect 372954 707398 373574 707482
rect 372954 707162 372986 707398
rect 373222 707162 373306 707398
rect 373542 707162 373574 707398
rect 372954 698614 373574 707162
rect 372954 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 373574 698614
rect 372954 698294 373574 698378
rect 372954 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 373574 698294
rect 372954 677977 373574 698058
rect 397794 704838 398414 711590
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 677977 398414 686898
rect 401514 705798 402134 711590
rect 401514 705562 401546 705798
rect 401782 705562 401866 705798
rect 402102 705562 402134 705798
rect 401514 705478 402134 705562
rect 401514 705242 401546 705478
rect 401782 705242 401866 705478
rect 402102 705242 402134 705478
rect 401514 691174 402134 705242
rect 401514 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 402134 691174
rect 401514 690854 402134 690938
rect 401514 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 402134 690854
rect 401514 677977 402134 690618
rect 405234 706758 405854 711590
rect 405234 706522 405266 706758
rect 405502 706522 405586 706758
rect 405822 706522 405854 706758
rect 405234 706438 405854 706522
rect 405234 706202 405266 706438
rect 405502 706202 405586 706438
rect 405822 706202 405854 706438
rect 405234 694894 405854 706202
rect 405234 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 405854 694894
rect 405234 694574 405854 694658
rect 405234 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 405854 694574
rect 405234 677977 405854 694338
rect 408954 707718 409574 711590
rect 408954 707482 408986 707718
rect 409222 707482 409306 707718
rect 409542 707482 409574 707718
rect 408954 707398 409574 707482
rect 408954 707162 408986 707398
rect 409222 707162 409306 707398
rect 409542 707162 409574 707398
rect 408954 698614 409574 707162
rect 408954 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 409574 698614
rect 408954 698294 409574 698378
rect 408954 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 409574 698294
rect 408954 677977 409574 698058
rect 433794 704838 434414 711590
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 677977 434414 686898
rect 437514 705798 438134 711590
rect 437514 705562 437546 705798
rect 437782 705562 437866 705798
rect 438102 705562 438134 705798
rect 437514 705478 438134 705562
rect 437514 705242 437546 705478
rect 437782 705242 437866 705478
rect 438102 705242 438134 705478
rect 437514 691174 438134 705242
rect 437514 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 438134 691174
rect 437514 690854 438134 690938
rect 437514 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 438134 690854
rect 437514 677977 438134 690618
rect 441234 706758 441854 711590
rect 441234 706522 441266 706758
rect 441502 706522 441586 706758
rect 441822 706522 441854 706758
rect 441234 706438 441854 706522
rect 441234 706202 441266 706438
rect 441502 706202 441586 706438
rect 441822 706202 441854 706438
rect 441234 694894 441854 706202
rect 441234 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 441854 694894
rect 441234 694574 441854 694658
rect 441234 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 441854 694574
rect 441234 677977 441854 694338
rect 444954 707718 445574 711590
rect 444954 707482 444986 707718
rect 445222 707482 445306 707718
rect 445542 707482 445574 707718
rect 444954 707398 445574 707482
rect 444954 707162 444986 707398
rect 445222 707162 445306 707398
rect 445542 707162 445574 707398
rect 444954 698614 445574 707162
rect 444954 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 445574 698614
rect 444954 698294 445574 698378
rect 444954 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 445574 698294
rect 444954 677977 445574 698058
rect 469794 704838 470414 711590
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 677977 470414 686898
rect 473514 705798 474134 711590
rect 473514 705562 473546 705798
rect 473782 705562 473866 705798
rect 474102 705562 474134 705798
rect 473514 705478 474134 705562
rect 473514 705242 473546 705478
rect 473782 705242 473866 705478
rect 474102 705242 474134 705478
rect 473514 691174 474134 705242
rect 473514 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 474134 691174
rect 473514 690854 474134 690938
rect 473514 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 474134 690854
rect 473514 677977 474134 690618
rect 477234 706758 477854 711590
rect 477234 706522 477266 706758
rect 477502 706522 477586 706758
rect 477822 706522 477854 706758
rect 477234 706438 477854 706522
rect 477234 706202 477266 706438
rect 477502 706202 477586 706438
rect 477822 706202 477854 706438
rect 477234 694894 477854 706202
rect 477234 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 477854 694894
rect 477234 694574 477854 694658
rect 477234 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 477854 694574
rect 477234 678332 477854 694338
rect 480954 707718 481574 711590
rect 480954 707482 480986 707718
rect 481222 707482 481306 707718
rect 481542 707482 481574 707718
rect 480954 707398 481574 707482
rect 480954 707162 480986 707398
rect 481222 707162 481306 707398
rect 481542 707162 481574 707398
rect 480954 698614 481574 707162
rect 480954 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 481574 698614
rect 480954 698294 481574 698378
rect 480954 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 481574 698294
rect 480954 677977 481574 698058
rect 505794 704838 506414 711590
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 677977 506414 686898
rect 509514 705798 510134 711590
rect 509514 705562 509546 705798
rect 509782 705562 509866 705798
rect 510102 705562 510134 705798
rect 509514 705478 510134 705562
rect 509514 705242 509546 705478
rect 509782 705242 509866 705478
rect 510102 705242 510134 705478
rect 509514 691174 510134 705242
rect 509514 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 510134 691174
rect 509514 690854 510134 690938
rect 509514 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 510134 690854
rect 509514 677977 510134 690618
rect 513234 706758 513854 711590
rect 513234 706522 513266 706758
rect 513502 706522 513586 706758
rect 513822 706522 513854 706758
rect 513234 706438 513854 706522
rect 513234 706202 513266 706438
rect 513502 706202 513586 706438
rect 513822 706202 513854 706438
rect 513234 694894 513854 706202
rect 513234 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 513854 694894
rect 513234 694574 513854 694658
rect 513234 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 513854 694574
rect 513234 677977 513854 694338
rect 516954 707718 517574 711590
rect 516954 707482 516986 707718
rect 517222 707482 517306 707718
rect 517542 707482 517574 707718
rect 516954 707398 517574 707482
rect 516954 707162 516986 707398
rect 517222 707162 517306 707398
rect 517542 707162 517574 707398
rect 516954 698614 517574 707162
rect 516954 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 517574 698614
rect 516954 698294 517574 698378
rect 516954 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 517574 698294
rect 516954 677977 517574 698058
rect 541794 704838 542414 711590
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 677977 542414 686898
rect 545514 705798 546134 711590
rect 545514 705562 545546 705798
rect 545782 705562 545866 705798
rect 546102 705562 546134 705798
rect 545514 705478 546134 705562
rect 545514 705242 545546 705478
rect 545782 705242 545866 705478
rect 546102 705242 546134 705478
rect 545514 691174 546134 705242
rect 545514 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 546134 691174
rect 545514 690854 546134 690938
rect 545514 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 546134 690854
rect 545514 677977 546134 690618
rect 549234 706758 549854 711590
rect 549234 706522 549266 706758
rect 549502 706522 549586 706758
rect 549822 706522 549854 706758
rect 549234 706438 549854 706522
rect 549234 706202 549266 706438
rect 549502 706202 549586 706438
rect 549822 706202 549854 706438
rect 549234 694894 549854 706202
rect 549234 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 549854 694894
rect 549234 694574 549854 694658
rect 549234 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 549854 694574
rect 549234 677977 549854 694338
rect 552954 707718 553574 711590
rect 552954 707482 552986 707718
rect 553222 707482 553306 707718
rect 553542 707482 553574 707718
rect 552954 707398 553574 707482
rect 552954 707162 552986 707398
rect 553222 707162 553306 707398
rect 553542 707162 553574 707398
rect 552954 698614 553574 707162
rect 552954 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 553574 698614
rect 552954 698294 553574 698378
rect 552954 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 553574 698294
rect 552954 677977 553574 698058
rect 567834 711558 568454 711590
rect 567834 711322 567866 711558
rect 568102 711322 568186 711558
rect 568422 711322 568454 711558
rect 567834 711238 568454 711322
rect 567834 711002 567866 711238
rect 568102 711002 568186 711238
rect 568422 711002 568454 711238
rect 9234 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 9854 658894
rect 9234 658574 9854 658658
rect 9234 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 9854 658574
rect 9234 622894 9854 658338
rect 567834 677494 568454 711002
rect 567834 677258 567866 677494
rect 568102 677258 568186 677494
rect 568422 677258 568454 677494
rect 567834 677174 568454 677258
rect 567834 676938 567866 677174
rect 568102 676938 568186 677174
rect 568422 676938 568454 677174
rect 31568 655174 31888 655206
rect 31568 654938 31610 655174
rect 31846 654938 31888 655174
rect 31568 654854 31888 654938
rect 31568 654618 31610 654854
rect 31846 654618 31888 654854
rect 31568 654586 31888 654618
rect 62288 655174 62608 655206
rect 62288 654938 62330 655174
rect 62566 654938 62608 655174
rect 62288 654854 62608 654938
rect 62288 654618 62330 654854
rect 62566 654618 62608 654854
rect 62288 654586 62608 654618
rect 93008 655174 93328 655206
rect 93008 654938 93050 655174
rect 93286 654938 93328 655174
rect 93008 654854 93328 654938
rect 93008 654618 93050 654854
rect 93286 654618 93328 654854
rect 93008 654586 93328 654618
rect 123728 655174 124048 655206
rect 123728 654938 123770 655174
rect 124006 654938 124048 655174
rect 123728 654854 124048 654938
rect 123728 654618 123770 654854
rect 124006 654618 124048 654854
rect 123728 654586 124048 654618
rect 154448 655174 154768 655206
rect 154448 654938 154490 655174
rect 154726 654938 154768 655174
rect 154448 654854 154768 654938
rect 154448 654618 154490 654854
rect 154726 654618 154768 654854
rect 154448 654586 154768 654618
rect 185168 655174 185488 655206
rect 185168 654938 185210 655174
rect 185446 654938 185488 655174
rect 185168 654854 185488 654938
rect 185168 654618 185210 654854
rect 185446 654618 185488 654854
rect 185168 654586 185488 654618
rect 215888 655174 216208 655206
rect 215888 654938 215930 655174
rect 216166 654938 216208 655174
rect 215888 654854 216208 654938
rect 215888 654618 215930 654854
rect 216166 654618 216208 654854
rect 215888 654586 216208 654618
rect 246608 655174 246928 655206
rect 246608 654938 246650 655174
rect 246886 654938 246928 655174
rect 246608 654854 246928 654938
rect 246608 654618 246650 654854
rect 246886 654618 246928 654854
rect 246608 654586 246928 654618
rect 277328 655174 277648 655206
rect 277328 654938 277370 655174
rect 277606 654938 277648 655174
rect 277328 654854 277648 654938
rect 277328 654618 277370 654854
rect 277606 654618 277648 654854
rect 277328 654586 277648 654618
rect 308048 655174 308368 655206
rect 308048 654938 308090 655174
rect 308326 654938 308368 655174
rect 308048 654854 308368 654938
rect 308048 654618 308090 654854
rect 308326 654618 308368 654854
rect 308048 654586 308368 654618
rect 338768 655174 339088 655206
rect 338768 654938 338810 655174
rect 339046 654938 339088 655174
rect 338768 654854 339088 654938
rect 338768 654618 338810 654854
rect 339046 654618 339088 654854
rect 338768 654586 339088 654618
rect 369488 655174 369808 655206
rect 369488 654938 369530 655174
rect 369766 654938 369808 655174
rect 369488 654854 369808 654938
rect 369488 654618 369530 654854
rect 369766 654618 369808 654854
rect 369488 654586 369808 654618
rect 400208 655174 400528 655206
rect 400208 654938 400250 655174
rect 400486 654938 400528 655174
rect 400208 654854 400528 654938
rect 400208 654618 400250 654854
rect 400486 654618 400528 654854
rect 400208 654586 400528 654618
rect 430928 655174 431248 655206
rect 430928 654938 430970 655174
rect 431206 654938 431248 655174
rect 430928 654854 431248 654938
rect 430928 654618 430970 654854
rect 431206 654618 431248 654854
rect 430928 654586 431248 654618
rect 461648 655174 461968 655206
rect 461648 654938 461690 655174
rect 461926 654938 461968 655174
rect 461648 654854 461968 654938
rect 461648 654618 461690 654854
rect 461926 654618 461968 654854
rect 461648 654586 461968 654618
rect 492368 655174 492688 655206
rect 492368 654938 492410 655174
rect 492646 654938 492688 655174
rect 492368 654854 492688 654938
rect 492368 654618 492410 654854
rect 492646 654618 492688 654854
rect 492368 654586 492688 654618
rect 523088 655174 523408 655206
rect 523088 654938 523130 655174
rect 523366 654938 523408 655174
rect 523088 654854 523408 654938
rect 523088 654618 523130 654854
rect 523366 654618 523408 654854
rect 523088 654586 523408 654618
rect 553808 655174 554128 655206
rect 553808 654938 553850 655174
rect 554086 654938 554128 655174
rect 553808 654854 554128 654938
rect 553808 654618 553850 654854
rect 554086 654618 554128 654854
rect 553808 654586 554128 654618
rect 16208 651454 16528 651486
rect 16208 651218 16250 651454
rect 16486 651218 16528 651454
rect 16208 651134 16528 651218
rect 16208 650898 16250 651134
rect 16486 650898 16528 651134
rect 16208 650866 16528 650898
rect 46928 651454 47248 651486
rect 46928 651218 46970 651454
rect 47206 651218 47248 651454
rect 46928 651134 47248 651218
rect 46928 650898 46970 651134
rect 47206 650898 47248 651134
rect 46928 650866 47248 650898
rect 77648 651454 77968 651486
rect 77648 651218 77690 651454
rect 77926 651218 77968 651454
rect 77648 651134 77968 651218
rect 77648 650898 77690 651134
rect 77926 650898 77968 651134
rect 77648 650866 77968 650898
rect 108368 651454 108688 651486
rect 108368 651218 108410 651454
rect 108646 651218 108688 651454
rect 108368 651134 108688 651218
rect 108368 650898 108410 651134
rect 108646 650898 108688 651134
rect 108368 650866 108688 650898
rect 139088 651454 139408 651486
rect 139088 651218 139130 651454
rect 139366 651218 139408 651454
rect 139088 651134 139408 651218
rect 139088 650898 139130 651134
rect 139366 650898 139408 651134
rect 139088 650866 139408 650898
rect 169808 651454 170128 651486
rect 169808 651218 169850 651454
rect 170086 651218 170128 651454
rect 169808 651134 170128 651218
rect 169808 650898 169850 651134
rect 170086 650898 170128 651134
rect 169808 650866 170128 650898
rect 200528 651454 200848 651486
rect 200528 651218 200570 651454
rect 200806 651218 200848 651454
rect 200528 651134 200848 651218
rect 200528 650898 200570 651134
rect 200806 650898 200848 651134
rect 200528 650866 200848 650898
rect 231248 651454 231568 651486
rect 231248 651218 231290 651454
rect 231526 651218 231568 651454
rect 231248 651134 231568 651218
rect 231248 650898 231290 651134
rect 231526 650898 231568 651134
rect 231248 650866 231568 650898
rect 261968 651454 262288 651486
rect 261968 651218 262010 651454
rect 262246 651218 262288 651454
rect 261968 651134 262288 651218
rect 261968 650898 262010 651134
rect 262246 650898 262288 651134
rect 261968 650866 262288 650898
rect 292688 651454 293008 651486
rect 292688 651218 292730 651454
rect 292966 651218 293008 651454
rect 292688 651134 293008 651218
rect 292688 650898 292730 651134
rect 292966 650898 293008 651134
rect 292688 650866 293008 650898
rect 323408 651454 323728 651486
rect 323408 651218 323450 651454
rect 323686 651218 323728 651454
rect 323408 651134 323728 651218
rect 323408 650898 323450 651134
rect 323686 650898 323728 651134
rect 323408 650866 323728 650898
rect 354128 651454 354448 651486
rect 354128 651218 354170 651454
rect 354406 651218 354448 651454
rect 354128 651134 354448 651218
rect 354128 650898 354170 651134
rect 354406 650898 354448 651134
rect 354128 650866 354448 650898
rect 384848 651454 385168 651486
rect 384848 651218 384890 651454
rect 385126 651218 385168 651454
rect 384848 651134 385168 651218
rect 384848 650898 384890 651134
rect 385126 650898 385168 651134
rect 384848 650866 385168 650898
rect 415568 651454 415888 651486
rect 415568 651218 415610 651454
rect 415846 651218 415888 651454
rect 415568 651134 415888 651218
rect 415568 650898 415610 651134
rect 415846 650898 415888 651134
rect 415568 650866 415888 650898
rect 446288 651454 446608 651486
rect 446288 651218 446330 651454
rect 446566 651218 446608 651454
rect 446288 651134 446608 651218
rect 446288 650898 446330 651134
rect 446566 650898 446608 651134
rect 446288 650866 446608 650898
rect 477008 651454 477328 651486
rect 477008 651218 477050 651454
rect 477286 651218 477328 651454
rect 477008 651134 477328 651218
rect 477008 650898 477050 651134
rect 477286 650898 477328 651134
rect 477008 650866 477328 650898
rect 507728 651454 508048 651486
rect 507728 651218 507770 651454
rect 508006 651218 508048 651454
rect 507728 651134 508048 651218
rect 507728 650898 507770 651134
rect 508006 650898 508048 651134
rect 507728 650866 508048 650898
rect 538448 651454 538768 651486
rect 538448 651218 538490 651454
rect 538726 651218 538768 651454
rect 538448 651134 538768 651218
rect 538448 650898 538490 651134
rect 538726 650898 538768 651134
rect 538448 650866 538768 650898
rect 9234 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 9854 622894
rect 9234 622574 9854 622658
rect 9234 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 9854 622574
rect 9234 586894 9854 622338
rect 567834 641494 568454 676938
rect 567834 641258 567866 641494
rect 568102 641258 568186 641494
rect 568422 641258 568454 641494
rect 567834 641174 568454 641258
rect 567834 640938 567866 641174
rect 568102 640938 568186 641174
rect 568422 640938 568454 641174
rect 31568 619174 31888 619206
rect 31568 618938 31610 619174
rect 31846 618938 31888 619174
rect 31568 618854 31888 618938
rect 31568 618618 31610 618854
rect 31846 618618 31888 618854
rect 31568 618586 31888 618618
rect 62288 619174 62608 619206
rect 62288 618938 62330 619174
rect 62566 618938 62608 619174
rect 62288 618854 62608 618938
rect 62288 618618 62330 618854
rect 62566 618618 62608 618854
rect 62288 618586 62608 618618
rect 93008 619174 93328 619206
rect 93008 618938 93050 619174
rect 93286 618938 93328 619174
rect 93008 618854 93328 618938
rect 93008 618618 93050 618854
rect 93286 618618 93328 618854
rect 93008 618586 93328 618618
rect 123728 619174 124048 619206
rect 123728 618938 123770 619174
rect 124006 618938 124048 619174
rect 123728 618854 124048 618938
rect 123728 618618 123770 618854
rect 124006 618618 124048 618854
rect 123728 618586 124048 618618
rect 154448 619174 154768 619206
rect 154448 618938 154490 619174
rect 154726 618938 154768 619174
rect 154448 618854 154768 618938
rect 154448 618618 154490 618854
rect 154726 618618 154768 618854
rect 154448 618586 154768 618618
rect 185168 619174 185488 619206
rect 185168 618938 185210 619174
rect 185446 618938 185488 619174
rect 185168 618854 185488 618938
rect 185168 618618 185210 618854
rect 185446 618618 185488 618854
rect 185168 618586 185488 618618
rect 215888 619174 216208 619206
rect 215888 618938 215930 619174
rect 216166 618938 216208 619174
rect 215888 618854 216208 618938
rect 215888 618618 215930 618854
rect 216166 618618 216208 618854
rect 215888 618586 216208 618618
rect 246608 619174 246928 619206
rect 246608 618938 246650 619174
rect 246886 618938 246928 619174
rect 246608 618854 246928 618938
rect 246608 618618 246650 618854
rect 246886 618618 246928 618854
rect 246608 618586 246928 618618
rect 277328 619174 277648 619206
rect 277328 618938 277370 619174
rect 277606 618938 277648 619174
rect 277328 618854 277648 618938
rect 277328 618618 277370 618854
rect 277606 618618 277648 618854
rect 277328 618586 277648 618618
rect 308048 619174 308368 619206
rect 308048 618938 308090 619174
rect 308326 618938 308368 619174
rect 308048 618854 308368 618938
rect 308048 618618 308090 618854
rect 308326 618618 308368 618854
rect 308048 618586 308368 618618
rect 338768 619174 339088 619206
rect 338768 618938 338810 619174
rect 339046 618938 339088 619174
rect 338768 618854 339088 618938
rect 338768 618618 338810 618854
rect 339046 618618 339088 618854
rect 338768 618586 339088 618618
rect 369488 619174 369808 619206
rect 369488 618938 369530 619174
rect 369766 618938 369808 619174
rect 369488 618854 369808 618938
rect 369488 618618 369530 618854
rect 369766 618618 369808 618854
rect 369488 618586 369808 618618
rect 400208 619174 400528 619206
rect 400208 618938 400250 619174
rect 400486 618938 400528 619174
rect 400208 618854 400528 618938
rect 400208 618618 400250 618854
rect 400486 618618 400528 618854
rect 400208 618586 400528 618618
rect 430928 619174 431248 619206
rect 430928 618938 430970 619174
rect 431206 618938 431248 619174
rect 430928 618854 431248 618938
rect 430928 618618 430970 618854
rect 431206 618618 431248 618854
rect 430928 618586 431248 618618
rect 461648 619174 461968 619206
rect 461648 618938 461690 619174
rect 461926 618938 461968 619174
rect 461648 618854 461968 618938
rect 461648 618618 461690 618854
rect 461926 618618 461968 618854
rect 461648 618586 461968 618618
rect 492368 619174 492688 619206
rect 492368 618938 492410 619174
rect 492646 618938 492688 619174
rect 492368 618854 492688 618938
rect 492368 618618 492410 618854
rect 492646 618618 492688 618854
rect 492368 618586 492688 618618
rect 523088 619174 523408 619206
rect 523088 618938 523130 619174
rect 523366 618938 523408 619174
rect 523088 618854 523408 618938
rect 523088 618618 523130 618854
rect 523366 618618 523408 618854
rect 523088 618586 523408 618618
rect 553808 619174 554128 619206
rect 553808 618938 553850 619174
rect 554086 618938 554128 619174
rect 553808 618854 554128 618938
rect 553808 618618 553850 618854
rect 554086 618618 554128 618854
rect 553808 618586 554128 618618
rect 16208 615454 16528 615486
rect 16208 615218 16250 615454
rect 16486 615218 16528 615454
rect 16208 615134 16528 615218
rect 16208 614898 16250 615134
rect 16486 614898 16528 615134
rect 16208 614866 16528 614898
rect 46928 615454 47248 615486
rect 46928 615218 46970 615454
rect 47206 615218 47248 615454
rect 46928 615134 47248 615218
rect 46928 614898 46970 615134
rect 47206 614898 47248 615134
rect 46928 614866 47248 614898
rect 77648 615454 77968 615486
rect 77648 615218 77690 615454
rect 77926 615218 77968 615454
rect 77648 615134 77968 615218
rect 77648 614898 77690 615134
rect 77926 614898 77968 615134
rect 77648 614866 77968 614898
rect 108368 615454 108688 615486
rect 108368 615218 108410 615454
rect 108646 615218 108688 615454
rect 108368 615134 108688 615218
rect 108368 614898 108410 615134
rect 108646 614898 108688 615134
rect 108368 614866 108688 614898
rect 139088 615454 139408 615486
rect 139088 615218 139130 615454
rect 139366 615218 139408 615454
rect 139088 615134 139408 615218
rect 139088 614898 139130 615134
rect 139366 614898 139408 615134
rect 139088 614866 139408 614898
rect 169808 615454 170128 615486
rect 169808 615218 169850 615454
rect 170086 615218 170128 615454
rect 169808 615134 170128 615218
rect 169808 614898 169850 615134
rect 170086 614898 170128 615134
rect 169808 614866 170128 614898
rect 200528 615454 200848 615486
rect 200528 615218 200570 615454
rect 200806 615218 200848 615454
rect 200528 615134 200848 615218
rect 200528 614898 200570 615134
rect 200806 614898 200848 615134
rect 200528 614866 200848 614898
rect 231248 615454 231568 615486
rect 231248 615218 231290 615454
rect 231526 615218 231568 615454
rect 231248 615134 231568 615218
rect 231248 614898 231290 615134
rect 231526 614898 231568 615134
rect 231248 614866 231568 614898
rect 261968 615454 262288 615486
rect 261968 615218 262010 615454
rect 262246 615218 262288 615454
rect 261968 615134 262288 615218
rect 261968 614898 262010 615134
rect 262246 614898 262288 615134
rect 261968 614866 262288 614898
rect 292688 615454 293008 615486
rect 292688 615218 292730 615454
rect 292966 615218 293008 615454
rect 292688 615134 293008 615218
rect 292688 614898 292730 615134
rect 292966 614898 293008 615134
rect 292688 614866 293008 614898
rect 323408 615454 323728 615486
rect 323408 615218 323450 615454
rect 323686 615218 323728 615454
rect 323408 615134 323728 615218
rect 323408 614898 323450 615134
rect 323686 614898 323728 615134
rect 323408 614866 323728 614898
rect 354128 615454 354448 615486
rect 354128 615218 354170 615454
rect 354406 615218 354448 615454
rect 354128 615134 354448 615218
rect 354128 614898 354170 615134
rect 354406 614898 354448 615134
rect 354128 614866 354448 614898
rect 384848 615454 385168 615486
rect 384848 615218 384890 615454
rect 385126 615218 385168 615454
rect 384848 615134 385168 615218
rect 384848 614898 384890 615134
rect 385126 614898 385168 615134
rect 384848 614866 385168 614898
rect 415568 615454 415888 615486
rect 415568 615218 415610 615454
rect 415846 615218 415888 615454
rect 415568 615134 415888 615218
rect 415568 614898 415610 615134
rect 415846 614898 415888 615134
rect 415568 614866 415888 614898
rect 446288 615454 446608 615486
rect 446288 615218 446330 615454
rect 446566 615218 446608 615454
rect 446288 615134 446608 615218
rect 446288 614898 446330 615134
rect 446566 614898 446608 615134
rect 446288 614866 446608 614898
rect 477008 615454 477328 615486
rect 477008 615218 477050 615454
rect 477286 615218 477328 615454
rect 477008 615134 477328 615218
rect 477008 614898 477050 615134
rect 477286 614898 477328 615134
rect 477008 614866 477328 614898
rect 507728 615454 508048 615486
rect 507728 615218 507770 615454
rect 508006 615218 508048 615454
rect 507728 615134 508048 615218
rect 507728 614898 507770 615134
rect 508006 614898 508048 615134
rect 507728 614866 508048 614898
rect 538448 615454 538768 615486
rect 538448 615218 538490 615454
rect 538726 615218 538768 615454
rect 538448 615134 538768 615218
rect 538448 614898 538490 615134
rect 538726 614898 538768 615134
rect 538448 614866 538768 614898
rect 9234 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 9854 586894
rect 9234 586574 9854 586658
rect 9234 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 9854 586574
rect 9234 550894 9854 586338
rect 567834 605494 568454 640938
rect 567834 605258 567866 605494
rect 568102 605258 568186 605494
rect 568422 605258 568454 605494
rect 567834 605174 568454 605258
rect 567834 604938 567866 605174
rect 568102 604938 568186 605174
rect 568422 604938 568454 605174
rect 31568 583174 31888 583206
rect 31568 582938 31610 583174
rect 31846 582938 31888 583174
rect 31568 582854 31888 582938
rect 31568 582618 31610 582854
rect 31846 582618 31888 582854
rect 31568 582586 31888 582618
rect 62288 583174 62608 583206
rect 62288 582938 62330 583174
rect 62566 582938 62608 583174
rect 62288 582854 62608 582938
rect 62288 582618 62330 582854
rect 62566 582618 62608 582854
rect 62288 582586 62608 582618
rect 93008 583174 93328 583206
rect 93008 582938 93050 583174
rect 93286 582938 93328 583174
rect 93008 582854 93328 582938
rect 93008 582618 93050 582854
rect 93286 582618 93328 582854
rect 93008 582586 93328 582618
rect 123728 583174 124048 583206
rect 123728 582938 123770 583174
rect 124006 582938 124048 583174
rect 123728 582854 124048 582938
rect 123728 582618 123770 582854
rect 124006 582618 124048 582854
rect 123728 582586 124048 582618
rect 154448 583174 154768 583206
rect 154448 582938 154490 583174
rect 154726 582938 154768 583174
rect 154448 582854 154768 582938
rect 154448 582618 154490 582854
rect 154726 582618 154768 582854
rect 154448 582586 154768 582618
rect 185168 583174 185488 583206
rect 185168 582938 185210 583174
rect 185446 582938 185488 583174
rect 185168 582854 185488 582938
rect 185168 582618 185210 582854
rect 185446 582618 185488 582854
rect 185168 582586 185488 582618
rect 215888 583174 216208 583206
rect 215888 582938 215930 583174
rect 216166 582938 216208 583174
rect 215888 582854 216208 582938
rect 215888 582618 215930 582854
rect 216166 582618 216208 582854
rect 215888 582586 216208 582618
rect 246608 583174 246928 583206
rect 246608 582938 246650 583174
rect 246886 582938 246928 583174
rect 246608 582854 246928 582938
rect 246608 582618 246650 582854
rect 246886 582618 246928 582854
rect 246608 582586 246928 582618
rect 277328 583174 277648 583206
rect 277328 582938 277370 583174
rect 277606 582938 277648 583174
rect 277328 582854 277648 582938
rect 277328 582618 277370 582854
rect 277606 582618 277648 582854
rect 277328 582586 277648 582618
rect 308048 583174 308368 583206
rect 308048 582938 308090 583174
rect 308326 582938 308368 583174
rect 308048 582854 308368 582938
rect 308048 582618 308090 582854
rect 308326 582618 308368 582854
rect 308048 582586 308368 582618
rect 338768 583174 339088 583206
rect 338768 582938 338810 583174
rect 339046 582938 339088 583174
rect 338768 582854 339088 582938
rect 338768 582618 338810 582854
rect 339046 582618 339088 582854
rect 338768 582586 339088 582618
rect 369488 583174 369808 583206
rect 369488 582938 369530 583174
rect 369766 582938 369808 583174
rect 369488 582854 369808 582938
rect 369488 582618 369530 582854
rect 369766 582618 369808 582854
rect 369488 582586 369808 582618
rect 400208 583174 400528 583206
rect 400208 582938 400250 583174
rect 400486 582938 400528 583174
rect 400208 582854 400528 582938
rect 400208 582618 400250 582854
rect 400486 582618 400528 582854
rect 400208 582586 400528 582618
rect 430928 583174 431248 583206
rect 430928 582938 430970 583174
rect 431206 582938 431248 583174
rect 430928 582854 431248 582938
rect 430928 582618 430970 582854
rect 431206 582618 431248 582854
rect 430928 582586 431248 582618
rect 461648 583174 461968 583206
rect 461648 582938 461690 583174
rect 461926 582938 461968 583174
rect 461648 582854 461968 582938
rect 461648 582618 461690 582854
rect 461926 582618 461968 582854
rect 461648 582586 461968 582618
rect 492368 583174 492688 583206
rect 492368 582938 492410 583174
rect 492646 582938 492688 583174
rect 492368 582854 492688 582938
rect 492368 582618 492410 582854
rect 492646 582618 492688 582854
rect 492368 582586 492688 582618
rect 523088 583174 523408 583206
rect 523088 582938 523130 583174
rect 523366 582938 523408 583174
rect 523088 582854 523408 582938
rect 523088 582618 523130 582854
rect 523366 582618 523408 582854
rect 523088 582586 523408 582618
rect 553808 583174 554128 583206
rect 553808 582938 553850 583174
rect 554086 582938 554128 583174
rect 553808 582854 554128 582938
rect 553808 582618 553850 582854
rect 554086 582618 554128 582854
rect 553808 582586 554128 582618
rect 16208 579454 16528 579486
rect 16208 579218 16250 579454
rect 16486 579218 16528 579454
rect 16208 579134 16528 579218
rect 16208 578898 16250 579134
rect 16486 578898 16528 579134
rect 16208 578866 16528 578898
rect 46928 579454 47248 579486
rect 46928 579218 46970 579454
rect 47206 579218 47248 579454
rect 46928 579134 47248 579218
rect 46928 578898 46970 579134
rect 47206 578898 47248 579134
rect 46928 578866 47248 578898
rect 77648 579454 77968 579486
rect 77648 579218 77690 579454
rect 77926 579218 77968 579454
rect 77648 579134 77968 579218
rect 77648 578898 77690 579134
rect 77926 578898 77968 579134
rect 77648 578866 77968 578898
rect 108368 579454 108688 579486
rect 108368 579218 108410 579454
rect 108646 579218 108688 579454
rect 108368 579134 108688 579218
rect 108368 578898 108410 579134
rect 108646 578898 108688 579134
rect 108368 578866 108688 578898
rect 139088 579454 139408 579486
rect 139088 579218 139130 579454
rect 139366 579218 139408 579454
rect 139088 579134 139408 579218
rect 139088 578898 139130 579134
rect 139366 578898 139408 579134
rect 139088 578866 139408 578898
rect 169808 579454 170128 579486
rect 169808 579218 169850 579454
rect 170086 579218 170128 579454
rect 169808 579134 170128 579218
rect 169808 578898 169850 579134
rect 170086 578898 170128 579134
rect 169808 578866 170128 578898
rect 200528 579454 200848 579486
rect 200528 579218 200570 579454
rect 200806 579218 200848 579454
rect 200528 579134 200848 579218
rect 200528 578898 200570 579134
rect 200806 578898 200848 579134
rect 200528 578866 200848 578898
rect 231248 579454 231568 579486
rect 231248 579218 231290 579454
rect 231526 579218 231568 579454
rect 231248 579134 231568 579218
rect 231248 578898 231290 579134
rect 231526 578898 231568 579134
rect 231248 578866 231568 578898
rect 261968 579454 262288 579486
rect 261968 579218 262010 579454
rect 262246 579218 262288 579454
rect 261968 579134 262288 579218
rect 261968 578898 262010 579134
rect 262246 578898 262288 579134
rect 261968 578866 262288 578898
rect 292688 579454 293008 579486
rect 292688 579218 292730 579454
rect 292966 579218 293008 579454
rect 292688 579134 293008 579218
rect 292688 578898 292730 579134
rect 292966 578898 293008 579134
rect 292688 578866 293008 578898
rect 323408 579454 323728 579486
rect 323408 579218 323450 579454
rect 323686 579218 323728 579454
rect 323408 579134 323728 579218
rect 323408 578898 323450 579134
rect 323686 578898 323728 579134
rect 323408 578866 323728 578898
rect 354128 579454 354448 579486
rect 354128 579218 354170 579454
rect 354406 579218 354448 579454
rect 354128 579134 354448 579218
rect 354128 578898 354170 579134
rect 354406 578898 354448 579134
rect 354128 578866 354448 578898
rect 384848 579454 385168 579486
rect 384848 579218 384890 579454
rect 385126 579218 385168 579454
rect 384848 579134 385168 579218
rect 384848 578898 384890 579134
rect 385126 578898 385168 579134
rect 384848 578866 385168 578898
rect 415568 579454 415888 579486
rect 415568 579218 415610 579454
rect 415846 579218 415888 579454
rect 415568 579134 415888 579218
rect 415568 578898 415610 579134
rect 415846 578898 415888 579134
rect 415568 578866 415888 578898
rect 446288 579454 446608 579486
rect 446288 579218 446330 579454
rect 446566 579218 446608 579454
rect 446288 579134 446608 579218
rect 446288 578898 446330 579134
rect 446566 578898 446608 579134
rect 446288 578866 446608 578898
rect 477008 579454 477328 579486
rect 477008 579218 477050 579454
rect 477286 579218 477328 579454
rect 477008 579134 477328 579218
rect 477008 578898 477050 579134
rect 477286 578898 477328 579134
rect 477008 578866 477328 578898
rect 507728 579454 508048 579486
rect 507728 579218 507770 579454
rect 508006 579218 508048 579454
rect 507728 579134 508048 579218
rect 507728 578898 507770 579134
rect 508006 578898 508048 579134
rect 507728 578866 508048 578898
rect 538448 579454 538768 579486
rect 538448 579218 538490 579454
rect 538726 579218 538768 579454
rect 538448 579134 538768 579218
rect 538448 578898 538490 579134
rect 538726 578898 538768 579134
rect 538448 578866 538768 578898
rect 9234 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 9854 550894
rect 9234 550574 9854 550658
rect 9234 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 9854 550574
rect 9234 514894 9854 550338
rect 567834 569494 568454 604938
rect 567834 569258 567866 569494
rect 568102 569258 568186 569494
rect 568422 569258 568454 569494
rect 567834 569174 568454 569258
rect 567834 568938 567866 569174
rect 568102 568938 568186 569174
rect 568422 568938 568454 569174
rect 31568 547174 31888 547206
rect 31568 546938 31610 547174
rect 31846 546938 31888 547174
rect 31568 546854 31888 546938
rect 31568 546618 31610 546854
rect 31846 546618 31888 546854
rect 31568 546586 31888 546618
rect 62288 547174 62608 547206
rect 62288 546938 62330 547174
rect 62566 546938 62608 547174
rect 62288 546854 62608 546938
rect 62288 546618 62330 546854
rect 62566 546618 62608 546854
rect 62288 546586 62608 546618
rect 93008 547174 93328 547206
rect 93008 546938 93050 547174
rect 93286 546938 93328 547174
rect 93008 546854 93328 546938
rect 93008 546618 93050 546854
rect 93286 546618 93328 546854
rect 93008 546586 93328 546618
rect 123728 547174 124048 547206
rect 123728 546938 123770 547174
rect 124006 546938 124048 547174
rect 123728 546854 124048 546938
rect 123728 546618 123770 546854
rect 124006 546618 124048 546854
rect 123728 546586 124048 546618
rect 154448 547174 154768 547206
rect 154448 546938 154490 547174
rect 154726 546938 154768 547174
rect 154448 546854 154768 546938
rect 154448 546618 154490 546854
rect 154726 546618 154768 546854
rect 154448 546586 154768 546618
rect 185168 547174 185488 547206
rect 185168 546938 185210 547174
rect 185446 546938 185488 547174
rect 185168 546854 185488 546938
rect 185168 546618 185210 546854
rect 185446 546618 185488 546854
rect 185168 546586 185488 546618
rect 215888 547174 216208 547206
rect 215888 546938 215930 547174
rect 216166 546938 216208 547174
rect 215888 546854 216208 546938
rect 215888 546618 215930 546854
rect 216166 546618 216208 546854
rect 215888 546586 216208 546618
rect 246608 547174 246928 547206
rect 246608 546938 246650 547174
rect 246886 546938 246928 547174
rect 246608 546854 246928 546938
rect 246608 546618 246650 546854
rect 246886 546618 246928 546854
rect 246608 546586 246928 546618
rect 277328 547174 277648 547206
rect 277328 546938 277370 547174
rect 277606 546938 277648 547174
rect 277328 546854 277648 546938
rect 277328 546618 277370 546854
rect 277606 546618 277648 546854
rect 277328 546586 277648 546618
rect 308048 547174 308368 547206
rect 308048 546938 308090 547174
rect 308326 546938 308368 547174
rect 308048 546854 308368 546938
rect 308048 546618 308090 546854
rect 308326 546618 308368 546854
rect 308048 546586 308368 546618
rect 338768 547174 339088 547206
rect 338768 546938 338810 547174
rect 339046 546938 339088 547174
rect 338768 546854 339088 546938
rect 338768 546618 338810 546854
rect 339046 546618 339088 546854
rect 338768 546586 339088 546618
rect 369488 547174 369808 547206
rect 369488 546938 369530 547174
rect 369766 546938 369808 547174
rect 369488 546854 369808 546938
rect 369488 546618 369530 546854
rect 369766 546618 369808 546854
rect 369488 546586 369808 546618
rect 400208 547174 400528 547206
rect 400208 546938 400250 547174
rect 400486 546938 400528 547174
rect 400208 546854 400528 546938
rect 400208 546618 400250 546854
rect 400486 546618 400528 546854
rect 400208 546586 400528 546618
rect 430928 547174 431248 547206
rect 430928 546938 430970 547174
rect 431206 546938 431248 547174
rect 430928 546854 431248 546938
rect 430928 546618 430970 546854
rect 431206 546618 431248 546854
rect 430928 546586 431248 546618
rect 461648 547174 461968 547206
rect 461648 546938 461690 547174
rect 461926 546938 461968 547174
rect 461648 546854 461968 546938
rect 461648 546618 461690 546854
rect 461926 546618 461968 546854
rect 461648 546586 461968 546618
rect 492368 547174 492688 547206
rect 492368 546938 492410 547174
rect 492646 546938 492688 547174
rect 492368 546854 492688 546938
rect 492368 546618 492410 546854
rect 492646 546618 492688 546854
rect 492368 546586 492688 546618
rect 523088 547174 523408 547206
rect 523088 546938 523130 547174
rect 523366 546938 523408 547174
rect 523088 546854 523408 546938
rect 523088 546618 523130 546854
rect 523366 546618 523408 546854
rect 523088 546586 523408 546618
rect 553808 547174 554128 547206
rect 553808 546938 553850 547174
rect 554086 546938 554128 547174
rect 553808 546854 554128 546938
rect 553808 546618 553850 546854
rect 554086 546618 554128 546854
rect 553808 546586 554128 546618
rect 16208 543454 16528 543486
rect 16208 543218 16250 543454
rect 16486 543218 16528 543454
rect 16208 543134 16528 543218
rect 16208 542898 16250 543134
rect 16486 542898 16528 543134
rect 16208 542866 16528 542898
rect 46928 543454 47248 543486
rect 46928 543218 46970 543454
rect 47206 543218 47248 543454
rect 46928 543134 47248 543218
rect 46928 542898 46970 543134
rect 47206 542898 47248 543134
rect 46928 542866 47248 542898
rect 77648 543454 77968 543486
rect 77648 543218 77690 543454
rect 77926 543218 77968 543454
rect 77648 543134 77968 543218
rect 77648 542898 77690 543134
rect 77926 542898 77968 543134
rect 77648 542866 77968 542898
rect 108368 543454 108688 543486
rect 108368 543218 108410 543454
rect 108646 543218 108688 543454
rect 108368 543134 108688 543218
rect 108368 542898 108410 543134
rect 108646 542898 108688 543134
rect 108368 542866 108688 542898
rect 139088 543454 139408 543486
rect 139088 543218 139130 543454
rect 139366 543218 139408 543454
rect 139088 543134 139408 543218
rect 139088 542898 139130 543134
rect 139366 542898 139408 543134
rect 139088 542866 139408 542898
rect 169808 543454 170128 543486
rect 169808 543218 169850 543454
rect 170086 543218 170128 543454
rect 169808 543134 170128 543218
rect 169808 542898 169850 543134
rect 170086 542898 170128 543134
rect 169808 542866 170128 542898
rect 200528 543454 200848 543486
rect 200528 543218 200570 543454
rect 200806 543218 200848 543454
rect 200528 543134 200848 543218
rect 200528 542898 200570 543134
rect 200806 542898 200848 543134
rect 200528 542866 200848 542898
rect 231248 543454 231568 543486
rect 231248 543218 231290 543454
rect 231526 543218 231568 543454
rect 231248 543134 231568 543218
rect 231248 542898 231290 543134
rect 231526 542898 231568 543134
rect 231248 542866 231568 542898
rect 261968 543454 262288 543486
rect 261968 543218 262010 543454
rect 262246 543218 262288 543454
rect 261968 543134 262288 543218
rect 261968 542898 262010 543134
rect 262246 542898 262288 543134
rect 261968 542866 262288 542898
rect 292688 543454 293008 543486
rect 292688 543218 292730 543454
rect 292966 543218 293008 543454
rect 292688 543134 293008 543218
rect 292688 542898 292730 543134
rect 292966 542898 293008 543134
rect 292688 542866 293008 542898
rect 323408 543454 323728 543486
rect 323408 543218 323450 543454
rect 323686 543218 323728 543454
rect 323408 543134 323728 543218
rect 323408 542898 323450 543134
rect 323686 542898 323728 543134
rect 323408 542866 323728 542898
rect 354128 543454 354448 543486
rect 354128 543218 354170 543454
rect 354406 543218 354448 543454
rect 354128 543134 354448 543218
rect 354128 542898 354170 543134
rect 354406 542898 354448 543134
rect 354128 542866 354448 542898
rect 384848 543454 385168 543486
rect 384848 543218 384890 543454
rect 385126 543218 385168 543454
rect 384848 543134 385168 543218
rect 384848 542898 384890 543134
rect 385126 542898 385168 543134
rect 384848 542866 385168 542898
rect 415568 543454 415888 543486
rect 415568 543218 415610 543454
rect 415846 543218 415888 543454
rect 415568 543134 415888 543218
rect 415568 542898 415610 543134
rect 415846 542898 415888 543134
rect 415568 542866 415888 542898
rect 446288 543454 446608 543486
rect 446288 543218 446330 543454
rect 446566 543218 446608 543454
rect 446288 543134 446608 543218
rect 446288 542898 446330 543134
rect 446566 542898 446608 543134
rect 446288 542866 446608 542898
rect 477008 543454 477328 543486
rect 477008 543218 477050 543454
rect 477286 543218 477328 543454
rect 477008 543134 477328 543218
rect 477008 542898 477050 543134
rect 477286 542898 477328 543134
rect 477008 542866 477328 542898
rect 507728 543454 508048 543486
rect 507728 543218 507770 543454
rect 508006 543218 508048 543454
rect 507728 543134 508048 543218
rect 507728 542898 507770 543134
rect 508006 542898 508048 543134
rect 507728 542866 508048 542898
rect 538448 543454 538768 543486
rect 538448 543218 538490 543454
rect 538726 543218 538768 543454
rect 538448 543134 538768 543218
rect 538448 542898 538490 543134
rect 538726 542898 538768 543134
rect 538448 542866 538768 542898
rect 9234 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 9854 514894
rect 9234 514574 9854 514658
rect 9234 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 9854 514574
rect 9234 478894 9854 514338
rect 567834 533494 568454 568938
rect 567834 533258 567866 533494
rect 568102 533258 568186 533494
rect 568422 533258 568454 533494
rect 567834 533174 568454 533258
rect 567834 532938 567866 533174
rect 568102 532938 568186 533174
rect 568422 532938 568454 533174
rect 31568 511174 31888 511206
rect 31568 510938 31610 511174
rect 31846 510938 31888 511174
rect 31568 510854 31888 510938
rect 31568 510618 31610 510854
rect 31846 510618 31888 510854
rect 31568 510586 31888 510618
rect 62288 511174 62608 511206
rect 62288 510938 62330 511174
rect 62566 510938 62608 511174
rect 62288 510854 62608 510938
rect 62288 510618 62330 510854
rect 62566 510618 62608 510854
rect 62288 510586 62608 510618
rect 93008 511174 93328 511206
rect 93008 510938 93050 511174
rect 93286 510938 93328 511174
rect 93008 510854 93328 510938
rect 93008 510618 93050 510854
rect 93286 510618 93328 510854
rect 93008 510586 93328 510618
rect 123728 511174 124048 511206
rect 123728 510938 123770 511174
rect 124006 510938 124048 511174
rect 123728 510854 124048 510938
rect 123728 510618 123770 510854
rect 124006 510618 124048 510854
rect 123728 510586 124048 510618
rect 154448 511174 154768 511206
rect 154448 510938 154490 511174
rect 154726 510938 154768 511174
rect 154448 510854 154768 510938
rect 154448 510618 154490 510854
rect 154726 510618 154768 510854
rect 154448 510586 154768 510618
rect 185168 511174 185488 511206
rect 185168 510938 185210 511174
rect 185446 510938 185488 511174
rect 185168 510854 185488 510938
rect 185168 510618 185210 510854
rect 185446 510618 185488 510854
rect 185168 510586 185488 510618
rect 215888 511174 216208 511206
rect 215888 510938 215930 511174
rect 216166 510938 216208 511174
rect 215888 510854 216208 510938
rect 215888 510618 215930 510854
rect 216166 510618 216208 510854
rect 215888 510586 216208 510618
rect 246608 511174 246928 511206
rect 246608 510938 246650 511174
rect 246886 510938 246928 511174
rect 246608 510854 246928 510938
rect 246608 510618 246650 510854
rect 246886 510618 246928 510854
rect 246608 510586 246928 510618
rect 277328 511174 277648 511206
rect 277328 510938 277370 511174
rect 277606 510938 277648 511174
rect 277328 510854 277648 510938
rect 277328 510618 277370 510854
rect 277606 510618 277648 510854
rect 277328 510586 277648 510618
rect 308048 511174 308368 511206
rect 308048 510938 308090 511174
rect 308326 510938 308368 511174
rect 308048 510854 308368 510938
rect 308048 510618 308090 510854
rect 308326 510618 308368 510854
rect 308048 510586 308368 510618
rect 338768 511174 339088 511206
rect 338768 510938 338810 511174
rect 339046 510938 339088 511174
rect 338768 510854 339088 510938
rect 338768 510618 338810 510854
rect 339046 510618 339088 510854
rect 338768 510586 339088 510618
rect 369488 511174 369808 511206
rect 369488 510938 369530 511174
rect 369766 510938 369808 511174
rect 369488 510854 369808 510938
rect 369488 510618 369530 510854
rect 369766 510618 369808 510854
rect 369488 510586 369808 510618
rect 400208 511174 400528 511206
rect 400208 510938 400250 511174
rect 400486 510938 400528 511174
rect 400208 510854 400528 510938
rect 400208 510618 400250 510854
rect 400486 510618 400528 510854
rect 400208 510586 400528 510618
rect 430928 511174 431248 511206
rect 430928 510938 430970 511174
rect 431206 510938 431248 511174
rect 430928 510854 431248 510938
rect 430928 510618 430970 510854
rect 431206 510618 431248 510854
rect 430928 510586 431248 510618
rect 461648 511174 461968 511206
rect 461648 510938 461690 511174
rect 461926 510938 461968 511174
rect 461648 510854 461968 510938
rect 461648 510618 461690 510854
rect 461926 510618 461968 510854
rect 461648 510586 461968 510618
rect 492368 511174 492688 511206
rect 492368 510938 492410 511174
rect 492646 510938 492688 511174
rect 492368 510854 492688 510938
rect 492368 510618 492410 510854
rect 492646 510618 492688 510854
rect 492368 510586 492688 510618
rect 523088 511174 523408 511206
rect 523088 510938 523130 511174
rect 523366 510938 523408 511174
rect 523088 510854 523408 510938
rect 523088 510618 523130 510854
rect 523366 510618 523408 510854
rect 523088 510586 523408 510618
rect 553808 511174 554128 511206
rect 553808 510938 553850 511174
rect 554086 510938 554128 511174
rect 553808 510854 554128 510938
rect 553808 510618 553850 510854
rect 554086 510618 554128 510854
rect 553808 510586 554128 510618
rect 16208 507454 16528 507486
rect 16208 507218 16250 507454
rect 16486 507218 16528 507454
rect 16208 507134 16528 507218
rect 16208 506898 16250 507134
rect 16486 506898 16528 507134
rect 16208 506866 16528 506898
rect 46928 507454 47248 507486
rect 46928 507218 46970 507454
rect 47206 507218 47248 507454
rect 46928 507134 47248 507218
rect 46928 506898 46970 507134
rect 47206 506898 47248 507134
rect 46928 506866 47248 506898
rect 77648 507454 77968 507486
rect 77648 507218 77690 507454
rect 77926 507218 77968 507454
rect 77648 507134 77968 507218
rect 77648 506898 77690 507134
rect 77926 506898 77968 507134
rect 77648 506866 77968 506898
rect 108368 507454 108688 507486
rect 108368 507218 108410 507454
rect 108646 507218 108688 507454
rect 108368 507134 108688 507218
rect 108368 506898 108410 507134
rect 108646 506898 108688 507134
rect 108368 506866 108688 506898
rect 139088 507454 139408 507486
rect 139088 507218 139130 507454
rect 139366 507218 139408 507454
rect 139088 507134 139408 507218
rect 139088 506898 139130 507134
rect 139366 506898 139408 507134
rect 139088 506866 139408 506898
rect 169808 507454 170128 507486
rect 169808 507218 169850 507454
rect 170086 507218 170128 507454
rect 169808 507134 170128 507218
rect 169808 506898 169850 507134
rect 170086 506898 170128 507134
rect 169808 506866 170128 506898
rect 200528 507454 200848 507486
rect 200528 507218 200570 507454
rect 200806 507218 200848 507454
rect 200528 507134 200848 507218
rect 200528 506898 200570 507134
rect 200806 506898 200848 507134
rect 200528 506866 200848 506898
rect 231248 507454 231568 507486
rect 231248 507218 231290 507454
rect 231526 507218 231568 507454
rect 231248 507134 231568 507218
rect 231248 506898 231290 507134
rect 231526 506898 231568 507134
rect 231248 506866 231568 506898
rect 261968 507454 262288 507486
rect 261968 507218 262010 507454
rect 262246 507218 262288 507454
rect 261968 507134 262288 507218
rect 261968 506898 262010 507134
rect 262246 506898 262288 507134
rect 261968 506866 262288 506898
rect 292688 507454 293008 507486
rect 292688 507218 292730 507454
rect 292966 507218 293008 507454
rect 292688 507134 293008 507218
rect 292688 506898 292730 507134
rect 292966 506898 293008 507134
rect 292688 506866 293008 506898
rect 323408 507454 323728 507486
rect 323408 507218 323450 507454
rect 323686 507218 323728 507454
rect 323408 507134 323728 507218
rect 323408 506898 323450 507134
rect 323686 506898 323728 507134
rect 323408 506866 323728 506898
rect 354128 507454 354448 507486
rect 354128 507218 354170 507454
rect 354406 507218 354448 507454
rect 354128 507134 354448 507218
rect 354128 506898 354170 507134
rect 354406 506898 354448 507134
rect 354128 506866 354448 506898
rect 384848 507454 385168 507486
rect 384848 507218 384890 507454
rect 385126 507218 385168 507454
rect 384848 507134 385168 507218
rect 384848 506898 384890 507134
rect 385126 506898 385168 507134
rect 384848 506866 385168 506898
rect 415568 507454 415888 507486
rect 415568 507218 415610 507454
rect 415846 507218 415888 507454
rect 415568 507134 415888 507218
rect 415568 506898 415610 507134
rect 415846 506898 415888 507134
rect 415568 506866 415888 506898
rect 446288 507454 446608 507486
rect 446288 507218 446330 507454
rect 446566 507218 446608 507454
rect 446288 507134 446608 507218
rect 446288 506898 446330 507134
rect 446566 506898 446608 507134
rect 446288 506866 446608 506898
rect 477008 507454 477328 507486
rect 477008 507218 477050 507454
rect 477286 507218 477328 507454
rect 477008 507134 477328 507218
rect 477008 506898 477050 507134
rect 477286 506898 477328 507134
rect 477008 506866 477328 506898
rect 507728 507454 508048 507486
rect 507728 507218 507770 507454
rect 508006 507218 508048 507454
rect 507728 507134 508048 507218
rect 507728 506898 507770 507134
rect 508006 506898 508048 507134
rect 507728 506866 508048 506898
rect 538448 507454 538768 507486
rect 538448 507218 538490 507454
rect 538726 507218 538768 507454
rect 538448 507134 538768 507218
rect 538448 506898 538490 507134
rect 538726 506898 538768 507134
rect 538448 506866 538768 506898
rect 9234 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 9854 478894
rect 9234 478574 9854 478658
rect 9234 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 9854 478574
rect 9234 442894 9854 478338
rect 567834 497494 568454 532938
rect 567834 497258 567866 497494
rect 568102 497258 568186 497494
rect 568422 497258 568454 497494
rect 567834 497174 568454 497258
rect 567834 496938 567866 497174
rect 568102 496938 568186 497174
rect 568422 496938 568454 497174
rect 31568 475174 31888 475206
rect 31568 474938 31610 475174
rect 31846 474938 31888 475174
rect 31568 474854 31888 474938
rect 31568 474618 31610 474854
rect 31846 474618 31888 474854
rect 31568 474586 31888 474618
rect 62288 475174 62608 475206
rect 62288 474938 62330 475174
rect 62566 474938 62608 475174
rect 62288 474854 62608 474938
rect 62288 474618 62330 474854
rect 62566 474618 62608 474854
rect 62288 474586 62608 474618
rect 93008 475174 93328 475206
rect 93008 474938 93050 475174
rect 93286 474938 93328 475174
rect 93008 474854 93328 474938
rect 93008 474618 93050 474854
rect 93286 474618 93328 474854
rect 93008 474586 93328 474618
rect 123728 475174 124048 475206
rect 123728 474938 123770 475174
rect 124006 474938 124048 475174
rect 123728 474854 124048 474938
rect 123728 474618 123770 474854
rect 124006 474618 124048 474854
rect 123728 474586 124048 474618
rect 154448 475174 154768 475206
rect 154448 474938 154490 475174
rect 154726 474938 154768 475174
rect 154448 474854 154768 474938
rect 154448 474618 154490 474854
rect 154726 474618 154768 474854
rect 154448 474586 154768 474618
rect 185168 475174 185488 475206
rect 185168 474938 185210 475174
rect 185446 474938 185488 475174
rect 185168 474854 185488 474938
rect 185168 474618 185210 474854
rect 185446 474618 185488 474854
rect 185168 474586 185488 474618
rect 215888 475174 216208 475206
rect 215888 474938 215930 475174
rect 216166 474938 216208 475174
rect 215888 474854 216208 474938
rect 215888 474618 215930 474854
rect 216166 474618 216208 474854
rect 215888 474586 216208 474618
rect 246608 475174 246928 475206
rect 246608 474938 246650 475174
rect 246886 474938 246928 475174
rect 246608 474854 246928 474938
rect 246608 474618 246650 474854
rect 246886 474618 246928 474854
rect 246608 474586 246928 474618
rect 277328 475174 277648 475206
rect 277328 474938 277370 475174
rect 277606 474938 277648 475174
rect 277328 474854 277648 474938
rect 277328 474618 277370 474854
rect 277606 474618 277648 474854
rect 277328 474586 277648 474618
rect 308048 475174 308368 475206
rect 308048 474938 308090 475174
rect 308326 474938 308368 475174
rect 308048 474854 308368 474938
rect 308048 474618 308090 474854
rect 308326 474618 308368 474854
rect 308048 474586 308368 474618
rect 338768 475174 339088 475206
rect 338768 474938 338810 475174
rect 339046 474938 339088 475174
rect 338768 474854 339088 474938
rect 338768 474618 338810 474854
rect 339046 474618 339088 474854
rect 338768 474586 339088 474618
rect 369488 475174 369808 475206
rect 369488 474938 369530 475174
rect 369766 474938 369808 475174
rect 369488 474854 369808 474938
rect 369488 474618 369530 474854
rect 369766 474618 369808 474854
rect 369488 474586 369808 474618
rect 400208 475174 400528 475206
rect 400208 474938 400250 475174
rect 400486 474938 400528 475174
rect 400208 474854 400528 474938
rect 400208 474618 400250 474854
rect 400486 474618 400528 474854
rect 400208 474586 400528 474618
rect 430928 475174 431248 475206
rect 430928 474938 430970 475174
rect 431206 474938 431248 475174
rect 430928 474854 431248 474938
rect 430928 474618 430970 474854
rect 431206 474618 431248 474854
rect 430928 474586 431248 474618
rect 461648 475174 461968 475206
rect 461648 474938 461690 475174
rect 461926 474938 461968 475174
rect 461648 474854 461968 474938
rect 461648 474618 461690 474854
rect 461926 474618 461968 474854
rect 461648 474586 461968 474618
rect 492368 475174 492688 475206
rect 492368 474938 492410 475174
rect 492646 474938 492688 475174
rect 492368 474854 492688 474938
rect 492368 474618 492410 474854
rect 492646 474618 492688 474854
rect 492368 474586 492688 474618
rect 523088 475174 523408 475206
rect 523088 474938 523130 475174
rect 523366 474938 523408 475174
rect 523088 474854 523408 474938
rect 523088 474618 523130 474854
rect 523366 474618 523408 474854
rect 523088 474586 523408 474618
rect 553808 475174 554128 475206
rect 553808 474938 553850 475174
rect 554086 474938 554128 475174
rect 553808 474854 554128 474938
rect 553808 474618 553850 474854
rect 554086 474618 554128 474854
rect 553808 474586 554128 474618
rect 16208 471454 16528 471486
rect 16208 471218 16250 471454
rect 16486 471218 16528 471454
rect 16208 471134 16528 471218
rect 16208 470898 16250 471134
rect 16486 470898 16528 471134
rect 16208 470866 16528 470898
rect 46928 471454 47248 471486
rect 46928 471218 46970 471454
rect 47206 471218 47248 471454
rect 46928 471134 47248 471218
rect 46928 470898 46970 471134
rect 47206 470898 47248 471134
rect 46928 470866 47248 470898
rect 77648 471454 77968 471486
rect 77648 471218 77690 471454
rect 77926 471218 77968 471454
rect 77648 471134 77968 471218
rect 77648 470898 77690 471134
rect 77926 470898 77968 471134
rect 77648 470866 77968 470898
rect 108368 471454 108688 471486
rect 108368 471218 108410 471454
rect 108646 471218 108688 471454
rect 108368 471134 108688 471218
rect 108368 470898 108410 471134
rect 108646 470898 108688 471134
rect 108368 470866 108688 470898
rect 139088 471454 139408 471486
rect 139088 471218 139130 471454
rect 139366 471218 139408 471454
rect 139088 471134 139408 471218
rect 139088 470898 139130 471134
rect 139366 470898 139408 471134
rect 139088 470866 139408 470898
rect 169808 471454 170128 471486
rect 169808 471218 169850 471454
rect 170086 471218 170128 471454
rect 169808 471134 170128 471218
rect 169808 470898 169850 471134
rect 170086 470898 170128 471134
rect 169808 470866 170128 470898
rect 200528 471454 200848 471486
rect 200528 471218 200570 471454
rect 200806 471218 200848 471454
rect 200528 471134 200848 471218
rect 200528 470898 200570 471134
rect 200806 470898 200848 471134
rect 200528 470866 200848 470898
rect 231248 471454 231568 471486
rect 231248 471218 231290 471454
rect 231526 471218 231568 471454
rect 231248 471134 231568 471218
rect 231248 470898 231290 471134
rect 231526 470898 231568 471134
rect 231248 470866 231568 470898
rect 261968 471454 262288 471486
rect 261968 471218 262010 471454
rect 262246 471218 262288 471454
rect 261968 471134 262288 471218
rect 261968 470898 262010 471134
rect 262246 470898 262288 471134
rect 261968 470866 262288 470898
rect 292688 471454 293008 471486
rect 292688 471218 292730 471454
rect 292966 471218 293008 471454
rect 292688 471134 293008 471218
rect 292688 470898 292730 471134
rect 292966 470898 293008 471134
rect 292688 470866 293008 470898
rect 323408 471454 323728 471486
rect 323408 471218 323450 471454
rect 323686 471218 323728 471454
rect 323408 471134 323728 471218
rect 323408 470898 323450 471134
rect 323686 470898 323728 471134
rect 323408 470866 323728 470898
rect 354128 471454 354448 471486
rect 354128 471218 354170 471454
rect 354406 471218 354448 471454
rect 354128 471134 354448 471218
rect 354128 470898 354170 471134
rect 354406 470898 354448 471134
rect 354128 470866 354448 470898
rect 384848 471454 385168 471486
rect 384848 471218 384890 471454
rect 385126 471218 385168 471454
rect 384848 471134 385168 471218
rect 384848 470898 384890 471134
rect 385126 470898 385168 471134
rect 384848 470866 385168 470898
rect 415568 471454 415888 471486
rect 415568 471218 415610 471454
rect 415846 471218 415888 471454
rect 415568 471134 415888 471218
rect 415568 470898 415610 471134
rect 415846 470898 415888 471134
rect 415568 470866 415888 470898
rect 446288 471454 446608 471486
rect 446288 471218 446330 471454
rect 446566 471218 446608 471454
rect 446288 471134 446608 471218
rect 446288 470898 446330 471134
rect 446566 470898 446608 471134
rect 446288 470866 446608 470898
rect 477008 471454 477328 471486
rect 477008 471218 477050 471454
rect 477286 471218 477328 471454
rect 477008 471134 477328 471218
rect 477008 470898 477050 471134
rect 477286 470898 477328 471134
rect 477008 470866 477328 470898
rect 507728 471454 508048 471486
rect 507728 471218 507770 471454
rect 508006 471218 508048 471454
rect 507728 471134 508048 471218
rect 507728 470898 507770 471134
rect 508006 470898 508048 471134
rect 507728 470866 508048 470898
rect 538448 471454 538768 471486
rect 538448 471218 538490 471454
rect 538726 471218 538768 471454
rect 538448 471134 538768 471218
rect 538448 470898 538490 471134
rect 538726 470898 538768 471134
rect 538448 470866 538768 470898
rect 9234 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 9854 442894
rect 9234 442574 9854 442658
rect 9234 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 9854 442574
rect 9234 406894 9854 442338
rect 567834 461494 568454 496938
rect 567834 461258 567866 461494
rect 568102 461258 568186 461494
rect 568422 461258 568454 461494
rect 567834 461174 568454 461258
rect 567834 460938 567866 461174
rect 568102 460938 568186 461174
rect 568422 460938 568454 461174
rect 31568 439174 31888 439206
rect 31568 438938 31610 439174
rect 31846 438938 31888 439174
rect 31568 438854 31888 438938
rect 31568 438618 31610 438854
rect 31846 438618 31888 438854
rect 31568 438586 31888 438618
rect 62288 439174 62608 439206
rect 62288 438938 62330 439174
rect 62566 438938 62608 439174
rect 62288 438854 62608 438938
rect 62288 438618 62330 438854
rect 62566 438618 62608 438854
rect 62288 438586 62608 438618
rect 93008 439174 93328 439206
rect 93008 438938 93050 439174
rect 93286 438938 93328 439174
rect 93008 438854 93328 438938
rect 93008 438618 93050 438854
rect 93286 438618 93328 438854
rect 93008 438586 93328 438618
rect 123728 439174 124048 439206
rect 123728 438938 123770 439174
rect 124006 438938 124048 439174
rect 123728 438854 124048 438938
rect 123728 438618 123770 438854
rect 124006 438618 124048 438854
rect 123728 438586 124048 438618
rect 154448 439174 154768 439206
rect 154448 438938 154490 439174
rect 154726 438938 154768 439174
rect 154448 438854 154768 438938
rect 154448 438618 154490 438854
rect 154726 438618 154768 438854
rect 154448 438586 154768 438618
rect 185168 439174 185488 439206
rect 185168 438938 185210 439174
rect 185446 438938 185488 439174
rect 185168 438854 185488 438938
rect 185168 438618 185210 438854
rect 185446 438618 185488 438854
rect 185168 438586 185488 438618
rect 215888 439174 216208 439206
rect 215888 438938 215930 439174
rect 216166 438938 216208 439174
rect 215888 438854 216208 438938
rect 215888 438618 215930 438854
rect 216166 438618 216208 438854
rect 215888 438586 216208 438618
rect 246608 439174 246928 439206
rect 246608 438938 246650 439174
rect 246886 438938 246928 439174
rect 246608 438854 246928 438938
rect 246608 438618 246650 438854
rect 246886 438618 246928 438854
rect 246608 438586 246928 438618
rect 277328 439174 277648 439206
rect 277328 438938 277370 439174
rect 277606 438938 277648 439174
rect 277328 438854 277648 438938
rect 277328 438618 277370 438854
rect 277606 438618 277648 438854
rect 277328 438586 277648 438618
rect 308048 439174 308368 439206
rect 308048 438938 308090 439174
rect 308326 438938 308368 439174
rect 308048 438854 308368 438938
rect 308048 438618 308090 438854
rect 308326 438618 308368 438854
rect 308048 438586 308368 438618
rect 338768 439174 339088 439206
rect 338768 438938 338810 439174
rect 339046 438938 339088 439174
rect 338768 438854 339088 438938
rect 338768 438618 338810 438854
rect 339046 438618 339088 438854
rect 338768 438586 339088 438618
rect 369488 439174 369808 439206
rect 369488 438938 369530 439174
rect 369766 438938 369808 439174
rect 369488 438854 369808 438938
rect 369488 438618 369530 438854
rect 369766 438618 369808 438854
rect 369488 438586 369808 438618
rect 400208 439174 400528 439206
rect 400208 438938 400250 439174
rect 400486 438938 400528 439174
rect 400208 438854 400528 438938
rect 400208 438618 400250 438854
rect 400486 438618 400528 438854
rect 400208 438586 400528 438618
rect 430928 439174 431248 439206
rect 430928 438938 430970 439174
rect 431206 438938 431248 439174
rect 430928 438854 431248 438938
rect 430928 438618 430970 438854
rect 431206 438618 431248 438854
rect 430928 438586 431248 438618
rect 461648 439174 461968 439206
rect 461648 438938 461690 439174
rect 461926 438938 461968 439174
rect 461648 438854 461968 438938
rect 461648 438618 461690 438854
rect 461926 438618 461968 438854
rect 461648 438586 461968 438618
rect 492368 439174 492688 439206
rect 492368 438938 492410 439174
rect 492646 438938 492688 439174
rect 492368 438854 492688 438938
rect 492368 438618 492410 438854
rect 492646 438618 492688 438854
rect 492368 438586 492688 438618
rect 523088 439174 523408 439206
rect 523088 438938 523130 439174
rect 523366 438938 523408 439174
rect 523088 438854 523408 438938
rect 523088 438618 523130 438854
rect 523366 438618 523408 438854
rect 523088 438586 523408 438618
rect 553808 439174 554128 439206
rect 553808 438938 553850 439174
rect 554086 438938 554128 439174
rect 553808 438854 554128 438938
rect 553808 438618 553850 438854
rect 554086 438618 554128 438854
rect 553808 438586 554128 438618
rect 16208 435454 16528 435486
rect 16208 435218 16250 435454
rect 16486 435218 16528 435454
rect 16208 435134 16528 435218
rect 16208 434898 16250 435134
rect 16486 434898 16528 435134
rect 16208 434866 16528 434898
rect 46928 435454 47248 435486
rect 46928 435218 46970 435454
rect 47206 435218 47248 435454
rect 46928 435134 47248 435218
rect 46928 434898 46970 435134
rect 47206 434898 47248 435134
rect 46928 434866 47248 434898
rect 77648 435454 77968 435486
rect 77648 435218 77690 435454
rect 77926 435218 77968 435454
rect 77648 435134 77968 435218
rect 77648 434898 77690 435134
rect 77926 434898 77968 435134
rect 77648 434866 77968 434898
rect 108368 435454 108688 435486
rect 108368 435218 108410 435454
rect 108646 435218 108688 435454
rect 108368 435134 108688 435218
rect 108368 434898 108410 435134
rect 108646 434898 108688 435134
rect 108368 434866 108688 434898
rect 139088 435454 139408 435486
rect 139088 435218 139130 435454
rect 139366 435218 139408 435454
rect 139088 435134 139408 435218
rect 139088 434898 139130 435134
rect 139366 434898 139408 435134
rect 139088 434866 139408 434898
rect 169808 435454 170128 435486
rect 169808 435218 169850 435454
rect 170086 435218 170128 435454
rect 169808 435134 170128 435218
rect 169808 434898 169850 435134
rect 170086 434898 170128 435134
rect 169808 434866 170128 434898
rect 200528 435454 200848 435486
rect 200528 435218 200570 435454
rect 200806 435218 200848 435454
rect 200528 435134 200848 435218
rect 200528 434898 200570 435134
rect 200806 434898 200848 435134
rect 200528 434866 200848 434898
rect 231248 435454 231568 435486
rect 231248 435218 231290 435454
rect 231526 435218 231568 435454
rect 231248 435134 231568 435218
rect 231248 434898 231290 435134
rect 231526 434898 231568 435134
rect 231248 434866 231568 434898
rect 261968 435454 262288 435486
rect 261968 435218 262010 435454
rect 262246 435218 262288 435454
rect 261968 435134 262288 435218
rect 261968 434898 262010 435134
rect 262246 434898 262288 435134
rect 261968 434866 262288 434898
rect 292688 435454 293008 435486
rect 292688 435218 292730 435454
rect 292966 435218 293008 435454
rect 292688 435134 293008 435218
rect 292688 434898 292730 435134
rect 292966 434898 293008 435134
rect 292688 434866 293008 434898
rect 323408 435454 323728 435486
rect 323408 435218 323450 435454
rect 323686 435218 323728 435454
rect 323408 435134 323728 435218
rect 323408 434898 323450 435134
rect 323686 434898 323728 435134
rect 323408 434866 323728 434898
rect 354128 435454 354448 435486
rect 354128 435218 354170 435454
rect 354406 435218 354448 435454
rect 354128 435134 354448 435218
rect 354128 434898 354170 435134
rect 354406 434898 354448 435134
rect 354128 434866 354448 434898
rect 384848 435454 385168 435486
rect 384848 435218 384890 435454
rect 385126 435218 385168 435454
rect 384848 435134 385168 435218
rect 384848 434898 384890 435134
rect 385126 434898 385168 435134
rect 384848 434866 385168 434898
rect 415568 435454 415888 435486
rect 415568 435218 415610 435454
rect 415846 435218 415888 435454
rect 415568 435134 415888 435218
rect 415568 434898 415610 435134
rect 415846 434898 415888 435134
rect 415568 434866 415888 434898
rect 446288 435454 446608 435486
rect 446288 435218 446330 435454
rect 446566 435218 446608 435454
rect 446288 435134 446608 435218
rect 446288 434898 446330 435134
rect 446566 434898 446608 435134
rect 446288 434866 446608 434898
rect 477008 435454 477328 435486
rect 477008 435218 477050 435454
rect 477286 435218 477328 435454
rect 477008 435134 477328 435218
rect 477008 434898 477050 435134
rect 477286 434898 477328 435134
rect 477008 434866 477328 434898
rect 507728 435454 508048 435486
rect 507728 435218 507770 435454
rect 508006 435218 508048 435454
rect 507728 435134 508048 435218
rect 507728 434898 507770 435134
rect 508006 434898 508048 435134
rect 507728 434866 508048 434898
rect 538448 435454 538768 435486
rect 538448 435218 538490 435454
rect 538726 435218 538768 435454
rect 538448 435134 538768 435218
rect 538448 434898 538490 435134
rect 538726 434898 538768 435134
rect 538448 434866 538768 434898
rect 9234 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 9854 406894
rect 9234 406574 9854 406658
rect 9234 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 9854 406574
rect 9234 370894 9854 406338
rect 567834 425494 568454 460938
rect 567834 425258 567866 425494
rect 568102 425258 568186 425494
rect 568422 425258 568454 425494
rect 567834 425174 568454 425258
rect 567834 424938 567866 425174
rect 568102 424938 568186 425174
rect 568422 424938 568454 425174
rect 31568 403174 31888 403206
rect 31568 402938 31610 403174
rect 31846 402938 31888 403174
rect 31568 402854 31888 402938
rect 31568 402618 31610 402854
rect 31846 402618 31888 402854
rect 31568 402586 31888 402618
rect 62288 403174 62608 403206
rect 62288 402938 62330 403174
rect 62566 402938 62608 403174
rect 62288 402854 62608 402938
rect 62288 402618 62330 402854
rect 62566 402618 62608 402854
rect 62288 402586 62608 402618
rect 93008 403174 93328 403206
rect 93008 402938 93050 403174
rect 93286 402938 93328 403174
rect 93008 402854 93328 402938
rect 93008 402618 93050 402854
rect 93286 402618 93328 402854
rect 93008 402586 93328 402618
rect 123728 403174 124048 403206
rect 123728 402938 123770 403174
rect 124006 402938 124048 403174
rect 123728 402854 124048 402938
rect 123728 402618 123770 402854
rect 124006 402618 124048 402854
rect 123728 402586 124048 402618
rect 154448 403174 154768 403206
rect 154448 402938 154490 403174
rect 154726 402938 154768 403174
rect 154448 402854 154768 402938
rect 154448 402618 154490 402854
rect 154726 402618 154768 402854
rect 154448 402586 154768 402618
rect 185168 403174 185488 403206
rect 185168 402938 185210 403174
rect 185446 402938 185488 403174
rect 185168 402854 185488 402938
rect 185168 402618 185210 402854
rect 185446 402618 185488 402854
rect 185168 402586 185488 402618
rect 215888 403174 216208 403206
rect 215888 402938 215930 403174
rect 216166 402938 216208 403174
rect 215888 402854 216208 402938
rect 215888 402618 215930 402854
rect 216166 402618 216208 402854
rect 215888 402586 216208 402618
rect 246608 403174 246928 403206
rect 246608 402938 246650 403174
rect 246886 402938 246928 403174
rect 246608 402854 246928 402938
rect 246608 402618 246650 402854
rect 246886 402618 246928 402854
rect 246608 402586 246928 402618
rect 277328 403174 277648 403206
rect 277328 402938 277370 403174
rect 277606 402938 277648 403174
rect 277328 402854 277648 402938
rect 277328 402618 277370 402854
rect 277606 402618 277648 402854
rect 277328 402586 277648 402618
rect 308048 403174 308368 403206
rect 308048 402938 308090 403174
rect 308326 402938 308368 403174
rect 308048 402854 308368 402938
rect 308048 402618 308090 402854
rect 308326 402618 308368 402854
rect 308048 402586 308368 402618
rect 338768 403174 339088 403206
rect 338768 402938 338810 403174
rect 339046 402938 339088 403174
rect 338768 402854 339088 402938
rect 338768 402618 338810 402854
rect 339046 402618 339088 402854
rect 338768 402586 339088 402618
rect 369488 403174 369808 403206
rect 369488 402938 369530 403174
rect 369766 402938 369808 403174
rect 369488 402854 369808 402938
rect 369488 402618 369530 402854
rect 369766 402618 369808 402854
rect 369488 402586 369808 402618
rect 400208 403174 400528 403206
rect 400208 402938 400250 403174
rect 400486 402938 400528 403174
rect 400208 402854 400528 402938
rect 400208 402618 400250 402854
rect 400486 402618 400528 402854
rect 400208 402586 400528 402618
rect 430928 403174 431248 403206
rect 430928 402938 430970 403174
rect 431206 402938 431248 403174
rect 430928 402854 431248 402938
rect 430928 402618 430970 402854
rect 431206 402618 431248 402854
rect 430928 402586 431248 402618
rect 461648 403174 461968 403206
rect 461648 402938 461690 403174
rect 461926 402938 461968 403174
rect 461648 402854 461968 402938
rect 461648 402618 461690 402854
rect 461926 402618 461968 402854
rect 461648 402586 461968 402618
rect 492368 403174 492688 403206
rect 492368 402938 492410 403174
rect 492646 402938 492688 403174
rect 492368 402854 492688 402938
rect 492368 402618 492410 402854
rect 492646 402618 492688 402854
rect 492368 402586 492688 402618
rect 523088 403174 523408 403206
rect 523088 402938 523130 403174
rect 523366 402938 523408 403174
rect 523088 402854 523408 402938
rect 523088 402618 523130 402854
rect 523366 402618 523408 402854
rect 523088 402586 523408 402618
rect 553808 403174 554128 403206
rect 553808 402938 553850 403174
rect 554086 402938 554128 403174
rect 553808 402854 554128 402938
rect 553808 402618 553850 402854
rect 554086 402618 554128 402854
rect 553808 402586 554128 402618
rect 16208 399454 16528 399486
rect 16208 399218 16250 399454
rect 16486 399218 16528 399454
rect 16208 399134 16528 399218
rect 16208 398898 16250 399134
rect 16486 398898 16528 399134
rect 16208 398866 16528 398898
rect 46928 399454 47248 399486
rect 46928 399218 46970 399454
rect 47206 399218 47248 399454
rect 46928 399134 47248 399218
rect 46928 398898 46970 399134
rect 47206 398898 47248 399134
rect 46928 398866 47248 398898
rect 77648 399454 77968 399486
rect 77648 399218 77690 399454
rect 77926 399218 77968 399454
rect 77648 399134 77968 399218
rect 77648 398898 77690 399134
rect 77926 398898 77968 399134
rect 77648 398866 77968 398898
rect 108368 399454 108688 399486
rect 108368 399218 108410 399454
rect 108646 399218 108688 399454
rect 108368 399134 108688 399218
rect 108368 398898 108410 399134
rect 108646 398898 108688 399134
rect 108368 398866 108688 398898
rect 139088 399454 139408 399486
rect 139088 399218 139130 399454
rect 139366 399218 139408 399454
rect 139088 399134 139408 399218
rect 139088 398898 139130 399134
rect 139366 398898 139408 399134
rect 139088 398866 139408 398898
rect 169808 399454 170128 399486
rect 169808 399218 169850 399454
rect 170086 399218 170128 399454
rect 169808 399134 170128 399218
rect 169808 398898 169850 399134
rect 170086 398898 170128 399134
rect 169808 398866 170128 398898
rect 200528 399454 200848 399486
rect 200528 399218 200570 399454
rect 200806 399218 200848 399454
rect 200528 399134 200848 399218
rect 200528 398898 200570 399134
rect 200806 398898 200848 399134
rect 200528 398866 200848 398898
rect 231248 399454 231568 399486
rect 231248 399218 231290 399454
rect 231526 399218 231568 399454
rect 231248 399134 231568 399218
rect 231248 398898 231290 399134
rect 231526 398898 231568 399134
rect 231248 398866 231568 398898
rect 261968 399454 262288 399486
rect 261968 399218 262010 399454
rect 262246 399218 262288 399454
rect 261968 399134 262288 399218
rect 261968 398898 262010 399134
rect 262246 398898 262288 399134
rect 261968 398866 262288 398898
rect 292688 399454 293008 399486
rect 292688 399218 292730 399454
rect 292966 399218 293008 399454
rect 292688 399134 293008 399218
rect 292688 398898 292730 399134
rect 292966 398898 293008 399134
rect 292688 398866 293008 398898
rect 323408 399454 323728 399486
rect 323408 399218 323450 399454
rect 323686 399218 323728 399454
rect 323408 399134 323728 399218
rect 323408 398898 323450 399134
rect 323686 398898 323728 399134
rect 323408 398866 323728 398898
rect 354128 399454 354448 399486
rect 354128 399218 354170 399454
rect 354406 399218 354448 399454
rect 354128 399134 354448 399218
rect 354128 398898 354170 399134
rect 354406 398898 354448 399134
rect 354128 398866 354448 398898
rect 384848 399454 385168 399486
rect 384848 399218 384890 399454
rect 385126 399218 385168 399454
rect 384848 399134 385168 399218
rect 384848 398898 384890 399134
rect 385126 398898 385168 399134
rect 384848 398866 385168 398898
rect 415568 399454 415888 399486
rect 415568 399218 415610 399454
rect 415846 399218 415888 399454
rect 415568 399134 415888 399218
rect 415568 398898 415610 399134
rect 415846 398898 415888 399134
rect 415568 398866 415888 398898
rect 446288 399454 446608 399486
rect 446288 399218 446330 399454
rect 446566 399218 446608 399454
rect 446288 399134 446608 399218
rect 446288 398898 446330 399134
rect 446566 398898 446608 399134
rect 446288 398866 446608 398898
rect 477008 399454 477328 399486
rect 477008 399218 477050 399454
rect 477286 399218 477328 399454
rect 477008 399134 477328 399218
rect 477008 398898 477050 399134
rect 477286 398898 477328 399134
rect 477008 398866 477328 398898
rect 507728 399454 508048 399486
rect 507728 399218 507770 399454
rect 508006 399218 508048 399454
rect 507728 399134 508048 399218
rect 507728 398898 507770 399134
rect 508006 398898 508048 399134
rect 507728 398866 508048 398898
rect 538448 399454 538768 399486
rect 538448 399218 538490 399454
rect 538726 399218 538768 399454
rect 538448 399134 538768 399218
rect 538448 398898 538490 399134
rect 538726 398898 538768 399134
rect 538448 398866 538768 398898
rect 9234 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 9854 370894
rect 9234 370574 9854 370658
rect 9234 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 9854 370574
rect 9234 334894 9854 370338
rect 567834 389494 568454 424938
rect 567834 389258 567866 389494
rect 568102 389258 568186 389494
rect 568422 389258 568454 389494
rect 567834 389174 568454 389258
rect 567834 388938 567866 389174
rect 568102 388938 568186 389174
rect 568422 388938 568454 389174
rect 31568 367174 31888 367206
rect 31568 366938 31610 367174
rect 31846 366938 31888 367174
rect 31568 366854 31888 366938
rect 31568 366618 31610 366854
rect 31846 366618 31888 366854
rect 31568 366586 31888 366618
rect 62288 367174 62608 367206
rect 62288 366938 62330 367174
rect 62566 366938 62608 367174
rect 62288 366854 62608 366938
rect 62288 366618 62330 366854
rect 62566 366618 62608 366854
rect 62288 366586 62608 366618
rect 93008 367174 93328 367206
rect 93008 366938 93050 367174
rect 93286 366938 93328 367174
rect 93008 366854 93328 366938
rect 93008 366618 93050 366854
rect 93286 366618 93328 366854
rect 93008 366586 93328 366618
rect 123728 367174 124048 367206
rect 123728 366938 123770 367174
rect 124006 366938 124048 367174
rect 123728 366854 124048 366938
rect 123728 366618 123770 366854
rect 124006 366618 124048 366854
rect 123728 366586 124048 366618
rect 154448 367174 154768 367206
rect 154448 366938 154490 367174
rect 154726 366938 154768 367174
rect 154448 366854 154768 366938
rect 154448 366618 154490 366854
rect 154726 366618 154768 366854
rect 154448 366586 154768 366618
rect 185168 367174 185488 367206
rect 185168 366938 185210 367174
rect 185446 366938 185488 367174
rect 185168 366854 185488 366938
rect 185168 366618 185210 366854
rect 185446 366618 185488 366854
rect 185168 366586 185488 366618
rect 215888 367174 216208 367206
rect 215888 366938 215930 367174
rect 216166 366938 216208 367174
rect 215888 366854 216208 366938
rect 215888 366618 215930 366854
rect 216166 366618 216208 366854
rect 215888 366586 216208 366618
rect 246608 367174 246928 367206
rect 246608 366938 246650 367174
rect 246886 366938 246928 367174
rect 246608 366854 246928 366938
rect 246608 366618 246650 366854
rect 246886 366618 246928 366854
rect 246608 366586 246928 366618
rect 277328 367174 277648 367206
rect 277328 366938 277370 367174
rect 277606 366938 277648 367174
rect 277328 366854 277648 366938
rect 277328 366618 277370 366854
rect 277606 366618 277648 366854
rect 277328 366586 277648 366618
rect 308048 367174 308368 367206
rect 308048 366938 308090 367174
rect 308326 366938 308368 367174
rect 308048 366854 308368 366938
rect 308048 366618 308090 366854
rect 308326 366618 308368 366854
rect 308048 366586 308368 366618
rect 338768 367174 339088 367206
rect 338768 366938 338810 367174
rect 339046 366938 339088 367174
rect 338768 366854 339088 366938
rect 338768 366618 338810 366854
rect 339046 366618 339088 366854
rect 338768 366586 339088 366618
rect 369488 367174 369808 367206
rect 369488 366938 369530 367174
rect 369766 366938 369808 367174
rect 369488 366854 369808 366938
rect 369488 366618 369530 366854
rect 369766 366618 369808 366854
rect 369488 366586 369808 366618
rect 400208 367174 400528 367206
rect 400208 366938 400250 367174
rect 400486 366938 400528 367174
rect 400208 366854 400528 366938
rect 400208 366618 400250 366854
rect 400486 366618 400528 366854
rect 400208 366586 400528 366618
rect 430928 367174 431248 367206
rect 430928 366938 430970 367174
rect 431206 366938 431248 367174
rect 430928 366854 431248 366938
rect 430928 366618 430970 366854
rect 431206 366618 431248 366854
rect 430928 366586 431248 366618
rect 461648 367174 461968 367206
rect 461648 366938 461690 367174
rect 461926 366938 461968 367174
rect 461648 366854 461968 366938
rect 461648 366618 461690 366854
rect 461926 366618 461968 366854
rect 461648 366586 461968 366618
rect 492368 367174 492688 367206
rect 492368 366938 492410 367174
rect 492646 366938 492688 367174
rect 492368 366854 492688 366938
rect 492368 366618 492410 366854
rect 492646 366618 492688 366854
rect 492368 366586 492688 366618
rect 523088 367174 523408 367206
rect 523088 366938 523130 367174
rect 523366 366938 523408 367174
rect 523088 366854 523408 366938
rect 523088 366618 523130 366854
rect 523366 366618 523408 366854
rect 523088 366586 523408 366618
rect 553808 367174 554128 367206
rect 553808 366938 553850 367174
rect 554086 366938 554128 367174
rect 553808 366854 554128 366938
rect 553808 366618 553850 366854
rect 554086 366618 554128 366854
rect 553808 366586 554128 366618
rect 16208 363454 16528 363486
rect 16208 363218 16250 363454
rect 16486 363218 16528 363454
rect 16208 363134 16528 363218
rect 16208 362898 16250 363134
rect 16486 362898 16528 363134
rect 16208 362866 16528 362898
rect 46928 363454 47248 363486
rect 46928 363218 46970 363454
rect 47206 363218 47248 363454
rect 46928 363134 47248 363218
rect 46928 362898 46970 363134
rect 47206 362898 47248 363134
rect 46928 362866 47248 362898
rect 77648 363454 77968 363486
rect 77648 363218 77690 363454
rect 77926 363218 77968 363454
rect 77648 363134 77968 363218
rect 77648 362898 77690 363134
rect 77926 362898 77968 363134
rect 77648 362866 77968 362898
rect 108368 363454 108688 363486
rect 108368 363218 108410 363454
rect 108646 363218 108688 363454
rect 108368 363134 108688 363218
rect 108368 362898 108410 363134
rect 108646 362898 108688 363134
rect 108368 362866 108688 362898
rect 139088 363454 139408 363486
rect 139088 363218 139130 363454
rect 139366 363218 139408 363454
rect 139088 363134 139408 363218
rect 139088 362898 139130 363134
rect 139366 362898 139408 363134
rect 139088 362866 139408 362898
rect 169808 363454 170128 363486
rect 169808 363218 169850 363454
rect 170086 363218 170128 363454
rect 169808 363134 170128 363218
rect 169808 362898 169850 363134
rect 170086 362898 170128 363134
rect 169808 362866 170128 362898
rect 200528 363454 200848 363486
rect 200528 363218 200570 363454
rect 200806 363218 200848 363454
rect 200528 363134 200848 363218
rect 200528 362898 200570 363134
rect 200806 362898 200848 363134
rect 200528 362866 200848 362898
rect 231248 363454 231568 363486
rect 231248 363218 231290 363454
rect 231526 363218 231568 363454
rect 231248 363134 231568 363218
rect 231248 362898 231290 363134
rect 231526 362898 231568 363134
rect 231248 362866 231568 362898
rect 261968 363454 262288 363486
rect 261968 363218 262010 363454
rect 262246 363218 262288 363454
rect 261968 363134 262288 363218
rect 261968 362898 262010 363134
rect 262246 362898 262288 363134
rect 261968 362866 262288 362898
rect 292688 363454 293008 363486
rect 292688 363218 292730 363454
rect 292966 363218 293008 363454
rect 292688 363134 293008 363218
rect 292688 362898 292730 363134
rect 292966 362898 293008 363134
rect 292688 362866 293008 362898
rect 323408 363454 323728 363486
rect 323408 363218 323450 363454
rect 323686 363218 323728 363454
rect 323408 363134 323728 363218
rect 323408 362898 323450 363134
rect 323686 362898 323728 363134
rect 323408 362866 323728 362898
rect 354128 363454 354448 363486
rect 354128 363218 354170 363454
rect 354406 363218 354448 363454
rect 354128 363134 354448 363218
rect 354128 362898 354170 363134
rect 354406 362898 354448 363134
rect 354128 362866 354448 362898
rect 384848 363454 385168 363486
rect 384848 363218 384890 363454
rect 385126 363218 385168 363454
rect 384848 363134 385168 363218
rect 384848 362898 384890 363134
rect 385126 362898 385168 363134
rect 384848 362866 385168 362898
rect 415568 363454 415888 363486
rect 415568 363218 415610 363454
rect 415846 363218 415888 363454
rect 415568 363134 415888 363218
rect 415568 362898 415610 363134
rect 415846 362898 415888 363134
rect 415568 362866 415888 362898
rect 446288 363454 446608 363486
rect 446288 363218 446330 363454
rect 446566 363218 446608 363454
rect 446288 363134 446608 363218
rect 446288 362898 446330 363134
rect 446566 362898 446608 363134
rect 446288 362866 446608 362898
rect 477008 363454 477328 363486
rect 477008 363218 477050 363454
rect 477286 363218 477328 363454
rect 477008 363134 477328 363218
rect 477008 362898 477050 363134
rect 477286 362898 477328 363134
rect 477008 362866 477328 362898
rect 507728 363454 508048 363486
rect 507728 363218 507770 363454
rect 508006 363218 508048 363454
rect 507728 363134 508048 363218
rect 507728 362898 507770 363134
rect 508006 362898 508048 363134
rect 507728 362866 508048 362898
rect 538448 363454 538768 363486
rect 538448 363218 538490 363454
rect 538726 363218 538768 363454
rect 538448 363134 538768 363218
rect 538448 362898 538490 363134
rect 538726 362898 538768 363134
rect 538448 362866 538768 362898
rect 9234 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 9854 334894
rect 9234 334574 9854 334658
rect 9234 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 9854 334574
rect 9234 298894 9854 334338
rect 567834 353494 568454 388938
rect 567834 353258 567866 353494
rect 568102 353258 568186 353494
rect 568422 353258 568454 353494
rect 567834 353174 568454 353258
rect 567834 352938 567866 353174
rect 568102 352938 568186 353174
rect 568422 352938 568454 353174
rect 31568 331174 31888 331206
rect 31568 330938 31610 331174
rect 31846 330938 31888 331174
rect 31568 330854 31888 330938
rect 31568 330618 31610 330854
rect 31846 330618 31888 330854
rect 31568 330586 31888 330618
rect 62288 331174 62608 331206
rect 62288 330938 62330 331174
rect 62566 330938 62608 331174
rect 62288 330854 62608 330938
rect 62288 330618 62330 330854
rect 62566 330618 62608 330854
rect 62288 330586 62608 330618
rect 93008 331174 93328 331206
rect 93008 330938 93050 331174
rect 93286 330938 93328 331174
rect 93008 330854 93328 330938
rect 93008 330618 93050 330854
rect 93286 330618 93328 330854
rect 93008 330586 93328 330618
rect 123728 331174 124048 331206
rect 123728 330938 123770 331174
rect 124006 330938 124048 331174
rect 123728 330854 124048 330938
rect 123728 330618 123770 330854
rect 124006 330618 124048 330854
rect 123728 330586 124048 330618
rect 154448 331174 154768 331206
rect 154448 330938 154490 331174
rect 154726 330938 154768 331174
rect 154448 330854 154768 330938
rect 154448 330618 154490 330854
rect 154726 330618 154768 330854
rect 154448 330586 154768 330618
rect 185168 331174 185488 331206
rect 185168 330938 185210 331174
rect 185446 330938 185488 331174
rect 185168 330854 185488 330938
rect 185168 330618 185210 330854
rect 185446 330618 185488 330854
rect 185168 330586 185488 330618
rect 215888 331174 216208 331206
rect 215888 330938 215930 331174
rect 216166 330938 216208 331174
rect 215888 330854 216208 330938
rect 215888 330618 215930 330854
rect 216166 330618 216208 330854
rect 215888 330586 216208 330618
rect 246608 331174 246928 331206
rect 246608 330938 246650 331174
rect 246886 330938 246928 331174
rect 246608 330854 246928 330938
rect 246608 330618 246650 330854
rect 246886 330618 246928 330854
rect 246608 330586 246928 330618
rect 277328 331174 277648 331206
rect 277328 330938 277370 331174
rect 277606 330938 277648 331174
rect 277328 330854 277648 330938
rect 277328 330618 277370 330854
rect 277606 330618 277648 330854
rect 277328 330586 277648 330618
rect 308048 331174 308368 331206
rect 308048 330938 308090 331174
rect 308326 330938 308368 331174
rect 308048 330854 308368 330938
rect 308048 330618 308090 330854
rect 308326 330618 308368 330854
rect 308048 330586 308368 330618
rect 338768 331174 339088 331206
rect 338768 330938 338810 331174
rect 339046 330938 339088 331174
rect 338768 330854 339088 330938
rect 338768 330618 338810 330854
rect 339046 330618 339088 330854
rect 338768 330586 339088 330618
rect 369488 331174 369808 331206
rect 369488 330938 369530 331174
rect 369766 330938 369808 331174
rect 369488 330854 369808 330938
rect 369488 330618 369530 330854
rect 369766 330618 369808 330854
rect 369488 330586 369808 330618
rect 400208 331174 400528 331206
rect 400208 330938 400250 331174
rect 400486 330938 400528 331174
rect 400208 330854 400528 330938
rect 400208 330618 400250 330854
rect 400486 330618 400528 330854
rect 400208 330586 400528 330618
rect 430928 331174 431248 331206
rect 430928 330938 430970 331174
rect 431206 330938 431248 331174
rect 430928 330854 431248 330938
rect 430928 330618 430970 330854
rect 431206 330618 431248 330854
rect 430928 330586 431248 330618
rect 461648 331174 461968 331206
rect 461648 330938 461690 331174
rect 461926 330938 461968 331174
rect 461648 330854 461968 330938
rect 461648 330618 461690 330854
rect 461926 330618 461968 330854
rect 461648 330586 461968 330618
rect 492368 331174 492688 331206
rect 492368 330938 492410 331174
rect 492646 330938 492688 331174
rect 492368 330854 492688 330938
rect 492368 330618 492410 330854
rect 492646 330618 492688 330854
rect 492368 330586 492688 330618
rect 523088 331174 523408 331206
rect 523088 330938 523130 331174
rect 523366 330938 523408 331174
rect 523088 330854 523408 330938
rect 523088 330618 523130 330854
rect 523366 330618 523408 330854
rect 523088 330586 523408 330618
rect 553808 331174 554128 331206
rect 553808 330938 553850 331174
rect 554086 330938 554128 331174
rect 553808 330854 554128 330938
rect 553808 330618 553850 330854
rect 554086 330618 554128 330854
rect 553808 330586 554128 330618
rect 16208 327454 16528 327486
rect 16208 327218 16250 327454
rect 16486 327218 16528 327454
rect 16208 327134 16528 327218
rect 16208 326898 16250 327134
rect 16486 326898 16528 327134
rect 16208 326866 16528 326898
rect 46928 327454 47248 327486
rect 46928 327218 46970 327454
rect 47206 327218 47248 327454
rect 46928 327134 47248 327218
rect 46928 326898 46970 327134
rect 47206 326898 47248 327134
rect 46928 326866 47248 326898
rect 77648 327454 77968 327486
rect 77648 327218 77690 327454
rect 77926 327218 77968 327454
rect 77648 327134 77968 327218
rect 77648 326898 77690 327134
rect 77926 326898 77968 327134
rect 77648 326866 77968 326898
rect 108368 327454 108688 327486
rect 108368 327218 108410 327454
rect 108646 327218 108688 327454
rect 108368 327134 108688 327218
rect 108368 326898 108410 327134
rect 108646 326898 108688 327134
rect 108368 326866 108688 326898
rect 139088 327454 139408 327486
rect 139088 327218 139130 327454
rect 139366 327218 139408 327454
rect 139088 327134 139408 327218
rect 139088 326898 139130 327134
rect 139366 326898 139408 327134
rect 139088 326866 139408 326898
rect 169808 327454 170128 327486
rect 169808 327218 169850 327454
rect 170086 327218 170128 327454
rect 169808 327134 170128 327218
rect 169808 326898 169850 327134
rect 170086 326898 170128 327134
rect 169808 326866 170128 326898
rect 200528 327454 200848 327486
rect 200528 327218 200570 327454
rect 200806 327218 200848 327454
rect 200528 327134 200848 327218
rect 200528 326898 200570 327134
rect 200806 326898 200848 327134
rect 200528 326866 200848 326898
rect 231248 327454 231568 327486
rect 231248 327218 231290 327454
rect 231526 327218 231568 327454
rect 231248 327134 231568 327218
rect 231248 326898 231290 327134
rect 231526 326898 231568 327134
rect 231248 326866 231568 326898
rect 261968 327454 262288 327486
rect 261968 327218 262010 327454
rect 262246 327218 262288 327454
rect 261968 327134 262288 327218
rect 261968 326898 262010 327134
rect 262246 326898 262288 327134
rect 261968 326866 262288 326898
rect 292688 327454 293008 327486
rect 292688 327218 292730 327454
rect 292966 327218 293008 327454
rect 292688 327134 293008 327218
rect 292688 326898 292730 327134
rect 292966 326898 293008 327134
rect 292688 326866 293008 326898
rect 323408 327454 323728 327486
rect 323408 327218 323450 327454
rect 323686 327218 323728 327454
rect 323408 327134 323728 327218
rect 323408 326898 323450 327134
rect 323686 326898 323728 327134
rect 323408 326866 323728 326898
rect 354128 327454 354448 327486
rect 354128 327218 354170 327454
rect 354406 327218 354448 327454
rect 354128 327134 354448 327218
rect 354128 326898 354170 327134
rect 354406 326898 354448 327134
rect 354128 326866 354448 326898
rect 384848 327454 385168 327486
rect 384848 327218 384890 327454
rect 385126 327218 385168 327454
rect 384848 327134 385168 327218
rect 384848 326898 384890 327134
rect 385126 326898 385168 327134
rect 384848 326866 385168 326898
rect 415568 327454 415888 327486
rect 415568 327218 415610 327454
rect 415846 327218 415888 327454
rect 415568 327134 415888 327218
rect 415568 326898 415610 327134
rect 415846 326898 415888 327134
rect 415568 326866 415888 326898
rect 446288 327454 446608 327486
rect 446288 327218 446330 327454
rect 446566 327218 446608 327454
rect 446288 327134 446608 327218
rect 446288 326898 446330 327134
rect 446566 326898 446608 327134
rect 446288 326866 446608 326898
rect 477008 327454 477328 327486
rect 477008 327218 477050 327454
rect 477286 327218 477328 327454
rect 477008 327134 477328 327218
rect 477008 326898 477050 327134
rect 477286 326898 477328 327134
rect 477008 326866 477328 326898
rect 507728 327454 508048 327486
rect 507728 327218 507770 327454
rect 508006 327218 508048 327454
rect 507728 327134 508048 327218
rect 507728 326898 507770 327134
rect 508006 326898 508048 327134
rect 507728 326866 508048 326898
rect 538448 327454 538768 327486
rect 538448 327218 538490 327454
rect 538726 327218 538768 327454
rect 538448 327134 538768 327218
rect 538448 326898 538490 327134
rect 538726 326898 538768 327134
rect 538448 326866 538768 326898
rect 9234 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 9854 298894
rect 9234 298574 9854 298658
rect 9234 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 9854 298574
rect 9234 262894 9854 298338
rect 567834 317494 568454 352938
rect 567834 317258 567866 317494
rect 568102 317258 568186 317494
rect 568422 317258 568454 317494
rect 567834 317174 568454 317258
rect 567834 316938 567866 317174
rect 568102 316938 568186 317174
rect 568422 316938 568454 317174
rect 31568 295174 31888 295206
rect 31568 294938 31610 295174
rect 31846 294938 31888 295174
rect 31568 294854 31888 294938
rect 31568 294618 31610 294854
rect 31846 294618 31888 294854
rect 31568 294586 31888 294618
rect 62288 295174 62608 295206
rect 62288 294938 62330 295174
rect 62566 294938 62608 295174
rect 62288 294854 62608 294938
rect 62288 294618 62330 294854
rect 62566 294618 62608 294854
rect 62288 294586 62608 294618
rect 93008 295174 93328 295206
rect 93008 294938 93050 295174
rect 93286 294938 93328 295174
rect 93008 294854 93328 294938
rect 93008 294618 93050 294854
rect 93286 294618 93328 294854
rect 93008 294586 93328 294618
rect 123728 295174 124048 295206
rect 123728 294938 123770 295174
rect 124006 294938 124048 295174
rect 123728 294854 124048 294938
rect 123728 294618 123770 294854
rect 124006 294618 124048 294854
rect 123728 294586 124048 294618
rect 154448 295174 154768 295206
rect 154448 294938 154490 295174
rect 154726 294938 154768 295174
rect 154448 294854 154768 294938
rect 154448 294618 154490 294854
rect 154726 294618 154768 294854
rect 154448 294586 154768 294618
rect 185168 295174 185488 295206
rect 185168 294938 185210 295174
rect 185446 294938 185488 295174
rect 185168 294854 185488 294938
rect 185168 294618 185210 294854
rect 185446 294618 185488 294854
rect 185168 294586 185488 294618
rect 215888 295174 216208 295206
rect 215888 294938 215930 295174
rect 216166 294938 216208 295174
rect 215888 294854 216208 294938
rect 215888 294618 215930 294854
rect 216166 294618 216208 294854
rect 215888 294586 216208 294618
rect 246608 295174 246928 295206
rect 246608 294938 246650 295174
rect 246886 294938 246928 295174
rect 246608 294854 246928 294938
rect 246608 294618 246650 294854
rect 246886 294618 246928 294854
rect 246608 294586 246928 294618
rect 277328 295174 277648 295206
rect 277328 294938 277370 295174
rect 277606 294938 277648 295174
rect 277328 294854 277648 294938
rect 277328 294618 277370 294854
rect 277606 294618 277648 294854
rect 277328 294586 277648 294618
rect 308048 295174 308368 295206
rect 308048 294938 308090 295174
rect 308326 294938 308368 295174
rect 308048 294854 308368 294938
rect 308048 294618 308090 294854
rect 308326 294618 308368 294854
rect 308048 294586 308368 294618
rect 338768 295174 339088 295206
rect 338768 294938 338810 295174
rect 339046 294938 339088 295174
rect 338768 294854 339088 294938
rect 338768 294618 338810 294854
rect 339046 294618 339088 294854
rect 338768 294586 339088 294618
rect 369488 295174 369808 295206
rect 369488 294938 369530 295174
rect 369766 294938 369808 295174
rect 369488 294854 369808 294938
rect 369488 294618 369530 294854
rect 369766 294618 369808 294854
rect 369488 294586 369808 294618
rect 400208 295174 400528 295206
rect 400208 294938 400250 295174
rect 400486 294938 400528 295174
rect 400208 294854 400528 294938
rect 400208 294618 400250 294854
rect 400486 294618 400528 294854
rect 400208 294586 400528 294618
rect 430928 295174 431248 295206
rect 430928 294938 430970 295174
rect 431206 294938 431248 295174
rect 430928 294854 431248 294938
rect 430928 294618 430970 294854
rect 431206 294618 431248 294854
rect 430928 294586 431248 294618
rect 461648 295174 461968 295206
rect 461648 294938 461690 295174
rect 461926 294938 461968 295174
rect 461648 294854 461968 294938
rect 461648 294618 461690 294854
rect 461926 294618 461968 294854
rect 461648 294586 461968 294618
rect 492368 295174 492688 295206
rect 492368 294938 492410 295174
rect 492646 294938 492688 295174
rect 492368 294854 492688 294938
rect 492368 294618 492410 294854
rect 492646 294618 492688 294854
rect 492368 294586 492688 294618
rect 523088 295174 523408 295206
rect 523088 294938 523130 295174
rect 523366 294938 523408 295174
rect 523088 294854 523408 294938
rect 523088 294618 523130 294854
rect 523366 294618 523408 294854
rect 523088 294586 523408 294618
rect 553808 295174 554128 295206
rect 553808 294938 553850 295174
rect 554086 294938 554128 295174
rect 553808 294854 554128 294938
rect 553808 294618 553850 294854
rect 554086 294618 554128 294854
rect 553808 294586 554128 294618
rect 16208 291454 16528 291486
rect 16208 291218 16250 291454
rect 16486 291218 16528 291454
rect 16208 291134 16528 291218
rect 16208 290898 16250 291134
rect 16486 290898 16528 291134
rect 16208 290866 16528 290898
rect 46928 291454 47248 291486
rect 46928 291218 46970 291454
rect 47206 291218 47248 291454
rect 46928 291134 47248 291218
rect 46928 290898 46970 291134
rect 47206 290898 47248 291134
rect 46928 290866 47248 290898
rect 77648 291454 77968 291486
rect 77648 291218 77690 291454
rect 77926 291218 77968 291454
rect 77648 291134 77968 291218
rect 77648 290898 77690 291134
rect 77926 290898 77968 291134
rect 77648 290866 77968 290898
rect 108368 291454 108688 291486
rect 108368 291218 108410 291454
rect 108646 291218 108688 291454
rect 108368 291134 108688 291218
rect 108368 290898 108410 291134
rect 108646 290898 108688 291134
rect 108368 290866 108688 290898
rect 139088 291454 139408 291486
rect 139088 291218 139130 291454
rect 139366 291218 139408 291454
rect 139088 291134 139408 291218
rect 139088 290898 139130 291134
rect 139366 290898 139408 291134
rect 139088 290866 139408 290898
rect 169808 291454 170128 291486
rect 169808 291218 169850 291454
rect 170086 291218 170128 291454
rect 169808 291134 170128 291218
rect 169808 290898 169850 291134
rect 170086 290898 170128 291134
rect 169808 290866 170128 290898
rect 200528 291454 200848 291486
rect 200528 291218 200570 291454
rect 200806 291218 200848 291454
rect 200528 291134 200848 291218
rect 200528 290898 200570 291134
rect 200806 290898 200848 291134
rect 200528 290866 200848 290898
rect 231248 291454 231568 291486
rect 231248 291218 231290 291454
rect 231526 291218 231568 291454
rect 231248 291134 231568 291218
rect 231248 290898 231290 291134
rect 231526 290898 231568 291134
rect 231248 290866 231568 290898
rect 261968 291454 262288 291486
rect 261968 291218 262010 291454
rect 262246 291218 262288 291454
rect 261968 291134 262288 291218
rect 261968 290898 262010 291134
rect 262246 290898 262288 291134
rect 261968 290866 262288 290898
rect 292688 291454 293008 291486
rect 292688 291218 292730 291454
rect 292966 291218 293008 291454
rect 292688 291134 293008 291218
rect 292688 290898 292730 291134
rect 292966 290898 293008 291134
rect 292688 290866 293008 290898
rect 323408 291454 323728 291486
rect 323408 291218 323450 291454
rect 323686 291218 323728 291454
rect 323408 291134 323728 291218
rect 323408 290898 323450 291134
rect 323686 290898 323728 291134
rect 323408 290866 323728 290898
rect 354128 291454 354448 291486
rect 354128 291218 354170 291454
rect 354406 291218 354448 291454
rect 354128 291134 354448 291218
rect 354128 290898 354170 291134
rect 354406 290898 354448 291134
rect 354128 290866 354448 290898
rect 384848 291454 385168 291486
rect 384848 291218 384890 291454
rect 385126 291218 385168 291454
rect 384848 291134 385168 291218
rect 384848 290898 384890 291134
rect 385126 290898 385168 291134
rect 384848 290866 385168 290898
rect 415568 291454 415888 291486
rect 415568 291218 415610 291454
rect 415846 291218 415888 291454
rect 415568 291134 415888 291218
rect 415568 290898 415610 291134
rect 415846 290898 415888 291134
rect 415568 290866 415888 290898
rect 446288 291454 446608 291486
rect 446288 291218 446330 291454
rect 446566 291218 446608 291454
rect 446288 291134 446608 291218
rect 446288 290898 446330 291134
rect 446566 290898 446608 291134
rect 446288 290866 446608 290898
rect 477008 291454 477328 291486
rect 477008 291218 477050 291454
rect 477286 291218 477328 291454
rect 477008 291134 477328 291218
rect 477008 290898 477050 291134
rect 477286 290898 477328 291134
rect 477008 290866 477328 290898
rect 507728 291454 508048 291486
rect 507728 291218 507770 291454
rect 508006 291218 508048 291454
rect 507728 291134 508048 291218
rect 507728 290898 507770 291134
rect 508006 290898 508048 291134
rect 507728 290866 508048 290898
rect 538448 291454 538768 291486
rect 538448 291218 538490 291454
rect 538726 291218 538768 291454
rect 538448 291134 538768 291218
rect 538448 290898 538490 291134
rect 538726 290898 538768 291134
rect 538448 290866 538768 290898
rect 9234 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 9854 262894
rect 9234 262574 9854 262658
rect 9234 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 9854 262574
rect 9234 226894 9854 262338
rect 567834 281494 568454 316938
rect 567834 281258 567866 281494
rect 568102 281258 568186 281494
rect 568422 281258 568454 281494
rect 567834 281174 568454 281258
rect 567834 280938 567866 281174
rect 568102 280938 568186 281174
rect 568422 280938 568454 281174
rect 31568 259174 31888 259206
rect 31568 258938 31610 259174
rect 31846 258938 31888 259174
rect 31568 258854 31888 258938
rect 31568 258618 31610 258854
rect 31846 258618 31888 258854
rect 31568 258586 31888 258618
rect 62288 259174 62608 259206
rect 62288 258938 62330 259174
rect 62566 258938 62608 259174
rect 62288 258854 62608 258938
rect 62288 258618 62330 258854
rect 62566 258618 62608 258854
rect 62288 258586 62608 258618
rect 93008 259174 93328 259206
rect 93008 258938 93050 259174
rect 93286 258938 93328 259174
rect 93008 258854 93328 258938
rect 93008 258618 93050 258854
rect 93286 258618 93328 258854
rect 93008 258586 93328 258618
rect 123728 259174 124048 259206
rect 123728 258938 123770 259174
rect 124006 258938 124048 259174
rect 123728 258854 124048 258938
rect 123728 258618 123770 258854
rect 124006 258618 124048 258854
rect 123728 258586 124048 258618
rect 154448 259174 154768 259206
rect 154448 258938 154490 259174
rect 154726 258938 154768 259174
rect 154448 258854 154768 258938
rect 154448 258618 154490 258854
rect 154726 258618 154768 258854
rect 154448 258586 154768 258618
rect 185168 259174 185488 259206
rect 185168 258938 185210 259174
rect 185446 258938 185488 259174
rect 185168 258854 185488 258938
rect 185168 258618 185210 258854
rect 185446 258618 185488 258854
rect 185168 258586 185488 258618
rect 215888 259174 216208 259206
rect 215888 258938 215930 259174
rect 216166 258938 216208 259174
rect 215888 258854 216208 258938
rect 215888 258618 215930 258854
rect 216166 258618 216208 258854
rect 215888 258586 216208 258618
rect 246608 259174 246928 259206
rect 246608 258938 246650 259174
rect 246886 258938 246928 259174
rect 246608 258854 246928 258938
rect 246608 258618 246650 258854
rect 246886 258618 246928 258854
rect 246608 258586 246928 258618
rect 277328 259174 277648 259206
rect 277328 258938 277370 259174
rect 277606 258938 277648 259174
rect 277328 258854 277648 258938
rect 277328 258618 277370 258854
rect 277606 258618 277648 258854
rect 277328 258586 277648 258618
rect 308048 259174 308368 259206
rect 308048 258938 308090 259174
rect 308326 258938 308368 259174
rect 308048 258854 308368 258938
rect 308048 258618 308090 258854
rect 308326 258618 308368 258854
rect 308048 258586 308368 258618
rect 338768 259174 339088 259206
rect 338768 258938 338810 259174
rect 339046 258938 339088 259174
rect 338768 258854 339088 258938
rect 338768 258618 338810 258854
rect 339046 258618 339088 258854
rect 338768 258586 339088 258618
rect 369488 259174 369808 259206
rect 369488 258938 369530 259174
rect 369766 258938 369808 259174
rect 369488 258854 369808 258938
rect 369488 258618 369530 258854
rect 369766 258618 369808 258854
rect 369488 258586 369808 258618
rect 400208 259174 400528 259206
rect 400208 258938 400250 259174
rect 400486 258938 400528 259174
rect 400208 258854 400528 258938
rect 400208 258618 400250 258854
rect 400486 258618 400528 258854
rect 400208 258586 400528 258618
rect 430928 259174 431248 259206
rect 430928 258938 430970 259174
rect 431206 258938 431248 259174
rect 430928 258854 431248 258938
rect 430928 258618 430970 258854
rect 431206 258618 431248 258854
rect 430928 258586 431248 258618
rect 461648 259174 461968 259206
rect 461648 258938 461690 259174
rect 461926 258938 461968 259174
rect 461648 258854 461968 258938
rect 461648 258618 461690 258854
rect 461926 258618 461968 258854
rect 461648 258586 461968 258618
rect 492368 259174 492688 259206
rect 492368 258938 492410 259174
rect 492646 258938 492688 259174
rect 492368 258854 492688 258938
rect 492368 258618 492410 258854
rect 492646 258618 492688 258854
rect 492368 258586 492688 258618
rect 523088 259174 523408 259206
rect 523088 258938 523130 259174
rect 523366 258938 523408 259174
rect 523088 258854 523408 258938
rect 523088 258618 523130 258854
rect 523366 258618 523408 258854
rect 523088 258586 523408 258618
rect 553808 259174 554128 259206
rect 553808 258938 553850 259174
rect 554086 258938 554128 259174
rect 553808 258854 554128 258938
rect 553808 258618 553850 258854
rect 554086 258618 554128 258854
rect 553808 258586 554128 258618
rect 16208 255454 16528 255486
rect 16208 255218 16250 255454
rect 16486 255218 16528 255454
rect 16208 255134 16528 255218
rect 16208 254898 16250 255134
rect 16486 254898 16528 255134
rect 16208 254866 16528 254898
rect 46928 255454 47248 255486
rect 46928 255218 46970 255454
rect 47206 255218 47248 255454
rect 46928 255134 47248 255218
rect 46928 254898 46970 255134
rect 47206 254898 47248 255134
rect 46928 254866 47248 254898
rect 77648 255454 77968 255486
rect 77648 255218 77690 255454
rect 77926 255218 77968 255454
rect 77648 255134 77968 255218
rect 77648 254898 77690 255134
rect 77926 254898 77968 255134
rect 77648 254866 77968 254898
rect 108368 255454 108688 255486
rect 108368 255218 108410 255454
rect 108646 255218 108688 255454
rect 108368 255134 108688 255218
rect 108368 254898 108410 255134
rect 108646 254898 108688 255134
rect 108368 254866 108688 254898
rect 139088 255454 139408 255486
rect 139088 255218 139130 255454
rect 139366 255218 139408 255454
rect 139088 255134 139408 255218
rect 139088 254898 139130 255134
rect 139366 254898 139408 255134
rect 139088 254866 139408 254898
rect 169808 255454 170128 255486
rect 169808 255218 169850 255454
rect 170086 255218 170128 255454
rect 169808 255134 170128 255218
rect 169808 254898 169850 255134
rect 170086 254898 170128 255134
rect 169808 254866 170128 254898
rect 200528 255454 200848 255486
rect 200528 255218 200570 255454
rect 200806 255218 200848 255454
rect 200528 255134 200848 255218
rect 200528 254898 200570 255134
rect 200806 254898 200848 255134
rect 200528 254866 200848 254898
rect 231248 255454 231568 255486
rect 231248 255218 231290 255454
rect 231526 255218 231568 255454
rect 231248 255134 231568 255218
rect 231248 254898 231290 255134
rect 231526 254898 231568 255134
rect 231248 254866 231568 254898
rect 261968 255454 262288 255486
rect 261968 255218 262010 255454
rect 262246 255218 262288 255454
rect 261968 255134 262288 255218
rect 261968 254898 262010 255134
rect 262246 254898 262288 255134
rect 261968 254866 262288 254898
rect 292688 255454 293008 255486
rect 292688 255218 292730 255454
rect 292966 255218 293008 255454
rect 292688 255134 293008 255218
rect 292688 254898 292730 255134
rect 292966 254898 293008 255134
rect 292688 254866 293008 254898
rect 323408 255454 323728 255486
rect 323408 255218 323450 255454
rect 323686 255218 323728 255454
rect 323408 255134 323728 255218
rect 323408 254898 323450 255134
rect 323686 254898 323728 255134
rect 323408 254866 323728 254898
rect 354128 255454 354448 255486
rect 354128 255218 354170 255454
rect 354406 255218 354448 255454
rect 354128 255134 354448 255218
rect 354128 254898 354170 255134
rect 354406 254898 354448 255134
rect 354128 254866 354448 254898
rect 384848 255454 385168 255486
rect 384848 255218 384890 255454
rect 385126 255218 385168 255454
rect 384848 255134 385168 255218
rect 384848 254898 384890 255134
rect 385126 254898 385168 255134
rect 384848 254866 385168 254898
rect 415568 255454 415888 255486
rect 415568 255218 415610 255454
rect 415846 255218 415888 255454
rect 415568 255134 415888 255218
rect 415568 254898 415610 255134
rect 415846 254898 415888 255134
rect 415568 254866 415888 254898
rect 446288 255454 446608 255486
rect 446288 255218 446330 255454
rect 446566 255218 446608 255454
rect 446288 255134 446608 255218
rect 446288 254898 446330 255134
rect 446566 254898 446608 255134
rect 446288 254866 446608 254898
rect 477008 255454 477328 255486
rect 477008 255218 477050 255454
rect 477286 255218 477328 255454
rect 477008 255134 477328 255218
rect 477008 254898 477050 255134
rect 477286 254898 477328 255134
rect 477008 254866 477328 254898
rect 507728 255454 508048 255486
rect 507728 255218 507770 255454
rect 508006 255218 508048 255454
rect 507728 255134 508048 255218
rect 507728 254898 507770 255134
rect 508006 254898 508048 255134
rect 507728 254866 508048 254898
rect 538448 255454 538768 255486
rect 538448 255218 538490 255454
rect 538726 255218 538768 255454
rect 538448 255134 538768 255218
rect 538448 254898 538490 255134
rect 538726 254898 538768 255134
rect 538448 254866 538768 254898
rect 9234 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 9854 226894
rect 9234 226574 9854 226658
rect 9234 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 9854 226574
rect 9234 190894 9854 226338
rect 567834 245494 568454 280938
rect 567834 245258 567866 245494
rect 568102 245258 568186 245494
rect 568422 245258 568454 245494
rect 567834 245174 568454 245258
rect 567834 244938 567866 245174
rect 568102 244938 568186 245174
rect 568422 244938 568454 245174
rect 31568 223174 31888 223206
rect 31568 222938 31610 223174
rect 31846 222938 31888 223174
rect 31568 222854 31888 222938
rect 31568 222618 31610 222854
rect 31846 222618 31888 222854
rect 31568 222586 31888 222618
rect 62288 223174 62608 223206
rect 62288 222938 62330 223174
rect 62566 222938 62608 223174
rect 62288 222854 62608 222938
rect 62288 222618 62330 222854
rect 62566 222618 62608 222854
rect 62288 222586 62608 222618
rect 93008 223174 93328 223206
rect 93008 222938 93050 223174
rect 93286 222938 93328 223174
rect 93008 222854 93328 222938
rect 93008 222618 93050 222854
rect 93286 222618 93328 222854
rect 93008 222586 93328 222618
rect 123728 223174 124048 223206
rect 123728 222938 123770 223174
rect 124006 222938 124048 223174
rect 123728 222854 124048 222938
rect 123728 222618 123770 222854
rect 124006 222618 124048 222854
rect 123728 222586 124048 222618
rect 154448 223174 154768 223206
rect 154448 222938 154490 223174
rect 154726 222938 154768 223174
rect 154448 222854 154768 222938
rect 154448 222618 154490 222854
rect 154726 222618 154768 222854
rect 154448 222586 154768 222618
rect 185168 223174 185488 223206
rect 185168 222938 185210 223174
rect 185446 222938 185488 223174
rect 185168 222854 185488 222938
rect 185168 222618 185210 222854
rect 185446 222618 185488 222854
rect 185168 222586 185488 222618
rect 215888 223174 216208 223206
rect 215888 222938 215930 223174
rect 216166 222938 216208 223174
rect 215888 222854 216208 222938
rect 215888 222618 215930 222854
rect 216166 222618 216208 222854
rect 215888 222586 216208 222618
rect 246608 223174 246928 223206
rect 246608 222938 246650 223174
rect 246886 222938 246928 223174
rect 246608 222854 246928 222938
rect 246608 222618 246650 222854
rect 246886 222618 246928 222854
rect 246608 222586 246928 222618
rect 277328 223174 277648 223206
rect 277328 222938 277370 223174
rect 277606 222938 277648 223174
rect 277328 222854 277648 222938
rect 277328 222618 277370 222854
rect 277606 222618 277648 222854
rect 277328 222586 277648 222618
rect 308048 223174 308368 223206
rect 308048 222938 308090 223174
rect 308326 222938 308368 223174
rect 308048 222854 308368 222938
rect 308048 222618 308090 222854
rect 308326 222618 308368 222854
rect 308048 222586 308368 222618
rect 338768 223174 339088 223206
rect 338768 222938 338810 223174
rect 339046 222938 339088 223174
rect 338768 222854 339088 222938
rect 338768 222618 338810 222854
rect 339046 222618 339088 222854
rect 338768 222586 339088 222618
rect 369488 223174 369808 223206
rect 369488 222938 369530 223174
rect 369766 222938 369808 223174
rect 369488 222854 369808 222938
rect 369488 222618 369530 222854
rect 369766 222618 369808 222854
rect 369488 222586 369808 222618
rect 400208 223174 400528 223206
rect 400208 222938 400250 223174
rect 400486 222938 400528 223174
rect 400208 222854 400528 222938
rect 400208 222618 400250 222854
rect 400486 222618 400528 222854
rect 400208 222586 400528 222618
rect 430928 223174 431248 223206
rect 430928 222938 430970 223174
rect 431206 222938 431248 223174
rect 430928 222854 431248 222938
rect 430928 222618 430970 222854
rect 431206 222618 431248 222854
rect 430928 222586 431248 222618
rect 461648 223174 461968 223206
rect 461648 222938 461690 223174
rect 461926 222938 461968 223174
rect 461648 222854 461968 222938
rect 461648 222618 461690 222854
rect 461926 222618 461968 222854
rect 461648 222586 461968 222618
rect 492368 223174 492688 223206
rect 492368 222938 492410 223174
rect 492646 222938 492688 223174
rect 492368 222854 492688 222938
rect 492368 222618 492410 222854
rect 492646 222618 492688 222854
rect 492368 222586 492688 222618
rect 523088 223174 523408 223206
rect 523088 222938 523130 223174
rect 523366 222938 523408 223174
rect 523088 222854 523408 222938
rect 523088 222618 523130 222854
rect 523366 222618 523408 222854
rect 523088 222586 523408 222618
rect 553808 223174 554128 223206
rect 553808 222938 553850 223174
rect 554086 222938 554128 223174
rect 553808 222854 554128 222938
rect 553808 222618 553850 222854
rect 554086 222618 554128 222854
rect 553808 222586 554128 222618
rect 16208 219454 16528 219486
rect 16208 219218 16250 219454
rect 16486 219218 16528 219454
rect 16208 219134 16528 219218
rect 16208 218898 16250 219134
rect 16486 218898 16528 219134
rect 16208 218866 16528 218898
rect 46928 219454 47248 219486
rect 46928 219218 46970 219454
rect 47206 219218 47248 219454
rect 46928 219134 47248 219218
rect 46928 218898 46970 219134
rect 47206 218898 47248 219134
rect 46928 218866 47248 218898
rect 77648 219454 77968 219486
rect 77648 219218 77690 219454
rect 77926 219218 77968 219454
rect 77648 219134 77968 219218
rect 77648 218898 77690 219134
rect 77926 218898 77968 219134
rect 77648 218866 77968 218898
rect 108368 219454 108688 219486
rect 108368 219218 108410 219454
rect 108646 219218 108688 219454
rect 108368 219134 108688 219218
rect 108368 218898 108410 219134
rect 108646 218898 108688 219134
rect 108368 218866 108688 218898
rect 139088 219454 139408 219486
rect 139088 219218 139130 219454
rect 139366 219218 139408 219454
rect 139088 219134 139408 219218
rect 139088 218898 139130 219134
rect 139366 218898 139408 219134
rect 139088 218866 139408 218898
rect 169808 219454 170128 219486
rect 169808 219218 169850 219454
rect 170086 219218 170128 219454
rect 169808 219134 170128 219218
rect 169808 218898 169850 219134
rect 170086 218898 170128 219134
rect 169808 218866 170128 218898
rect 200528 219454 200848 219486
rect 200528 219218 200570 219454
rect 200806 219218 200848 219454
rect 200528 219134 200848 219218
rect 200528 218898 200570 219134
rect 200806 218898 200848 219134
rect 200528 218866 200848 218898
rect 231248 219454 231568 219486
rect 231248 219218 231290 219454
rect 231526 219218 231568 219454
rect 231248 219134 231568 219218
rect 231248 218898 231290 219134
rect 231526 218898 231568 219134
rect 231248 218866 231568 218898
rect 261968 219454 262288 219486
rect 261968 219218 262010 219454
rect 262246 219218 262288 219454
rect 261968 219134 262288 219218
rect 261968 218898 262010 219134
rect 262246 218898 262288 219134
rect 261968 218866 262288 218898
rect 292688 219454 293008 219486
rect 292688 219218 292730 219454
rect 292966 219218 293008 219454
rect 292688 219134 293008 219218
rect 292688 218898 292730 219134
rect 292966 218898 293008 219134
rect 292688 218866 293008 218898
rect 323408 219454 323728 219486
rect 323408 219218 323450 219454
rect 323686 219218 323728 219454
rect 323408 219134 323728 219218
rect 323408 218898 323450 219134
rect 323686 218898 323728 219134
rect 323408 218866 323728 218898
rect 354128 219454 354448 219486
rect 354128 219218 354170 219454
rect 354406 219218 354448 219454
rect 354128 219134 354448 219218
rect 354128 218898 354170 219134
rect 354406 218898 354448 219134
rect 354128 218866 354448 218898
rect 384848 219454 385168 219486
rect 384848 219218 384890 219454
rect 385126 219218 385168 219454
rect 384848 219134 385168 219218
rect 384848 218898 384890 219134
rect 385126 218898 385168 219134
rect 384848 218866 385168 218898
rect 415568 219454 415888 219486
rect 415568 219218 415610 219454
rect 415846 219218 415888 219454
rect 415568 219134 415888 219218
rect 415568 218898 415610 219134
rect 415846 218898 415888 219134
rect 415568 218866 415888 218898
rect 446288 219454 446608 219486
rect 446288 219218 446330 219454
rect 446566 219218 446608 219454
rect 446288 219134 446608 219218
rect 446288 218898 446330 219134
rect 446566 218898 446608 219134
rect 446288 218866 446608 218898
rect 477008 219454 477328 219486
rect 477008 219218 477050 219454
rect 477286 219218 477328 219454
rect 477008 219134 477328 219218
rect 477008 218898 477050 219134
rect 477286 218898 477328 219134
rect 477008 218866 477328 218898
rect 507728 219454 508048 219486
rect 507728 219218 507770 219454
rect 508006 219218 508048 219454
rect 507728 219134 508048 219218
rect 507728 218898 507770 219134
rect 508006 218898 508048 219134
rect 507728 218866 508048 218898
rect 538448 219454 538768 219486
rect 538448 219218 538490 219454
rect 538726 219218 538768 219454
rect 538448 219134 538768 219218
rect 538448 218898 538490 219134
rect 538726 218898 538768 219134
rect 538448 218866 538768 218898
rect 9234 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 9854 190894
rect 9234 190574 9854 190658
rect 9234 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 9854 190574
rect 9234 154894 9854 190338
rect 567834 209494 568454 244938
rect 567834 209258 567866 209494
rect 568102 209258 568186 209494
rect 568422 209258 568454 209494
rect 567834 209174 568454 209258
rect 567834 208938 567866 209174
rect 568102 208938 568186 209174
rect 568422 208938 568454 209174
rect 31568 187174 31888 187206
rect 31568 186938 31610 187174
rect 31846 186938 31888 187174
rect 31568 186854 31888 186938
rect 31568 186618 31610 186854
rect 31846 186618 31888 186854
rect 31568 186586 31888 186618
rect 62288 187174 62608 187206
rect 62288 186938 62330 187174
rect 62566 186938 62608 187174
rect 62288 186854 62608 186938
rect 62288 186618 62330 186854
rect 62566 186618 62608 186854
rect 62288 186586 62608 186618
rect 93008 187174 93328 187206
rect 93008 186938 93050 187174
rect 93286 186938 93328 187174
rect 93008 186854 93328 186938
rect 93008 186618 93050 186854
rect 93286 186618 93328 186854
rect 93008 186586 93328 186618
rect 123728 187174 124048 187206
rect 123728 186938 123770 187174
rect 124006 186938 124048 187174
rect 123728 186854 124048 186938
rect 123728 186618 123770 186854
rect 124006 186618 124048 186854
rect 123728 186586 124048 186618
rect 154448 187174 154768 187206
rect 154448 186938 154490 187174
rect 154726 186938 154768 187174
rect 154448 186854 154768 186938
rect 154448 186618 154490 186854
rect 154726 186618 154768 186854
rect 154448 186586 154768 186618
rect 185168 187174 185488 187206
rect 185168 186938 185210 187174
rect 185446 186938 185488 187174
rect 185168 186854 185488 186938
rect 185168 186618 185210 186854
rect 185446 186618 185488 186854
rect 185168 186586 185488 186618
rect 215888 187174 216208 187206
rect 215888 186938 215930 187174
rect 216166 186938 216208 187174
rect 215888 186854 216208 186938
rect 215888 186618 215930 186854
rect 216166 186618 216208 186854
rect 215888 186586 216208 186618
rect 246608 187174 246928 187206
rect 246608 186938 246650 187174
rect 246886 186938 246928 187174
rect 246608 186854 246928 186938
rect 246608 186618 246650 186854
rect 246886 186618 246928 186854
rect 246608 186586 246928 186618
rect 277328 187174 277648 187206
rect 277328 186938 277370 187174
rect 277606 186938 277648 187174
rect 277328 186854 277648 186938
rect 277328 186618 277370 186854
rect 277606 186618 277648 186854
rect 277328 186586 277648 186618
rect 308048 187174 308368 187206
rect 308048 186938 308090 187174
rect 308326 186938 308368 187174
rect 308048 186854 308368 186938
rect 308048 186618 308090 186854
rect 308326 186618 308368 186854
rect 308048 186586 308368 186618
rect 338768 187174 339088 187206
rect 338768 186938 338810 187174
rect 339046 186938 339088 187174
rect 338768 186854 339088 186938
rect 338768 186618 338810 186854
rect 339046 186618 339088 186854
rect 338768 186586 339088 186618
rect 369488 187174 369808 187206
rect 369488 186938 369530 187174
rect 369766 186938 369808 187174
rect 369488 186854 369808 186938
rect 369488 186618 369530 186854
rect 369766 186618 369808 186854
rect 369488 186586 369808 186618
rect 400208 187174 400528 187206
rect 400208 186938 400250 187174
rect 400486 186938 400528 187174
rect 400208 186854 400528 186938
rect 400208 186618 400250 186854
rect 400486 186618 400528 186854
rect 400208 186586 400528 186618
rect 430928 187174 431248 187206
rect 430928 186938 430970 187174
rect 431206 186938 431248 187174
rect 430928 186854 431248 186938
rect 430928 186618 430970 186854
rect 431206 186618 431248 186854
rect 430928 186586 431248 186618
rect 461648 187174 461968 187206
rect 461648 186938 461690 187174
rect 461926 186938 461968 187174
rect 461648 186854 461968 186938
rect 461648 186618 461690 186854
rect 461926 186618 461968 186854
rect 461648 186586 461968 186618
rect 492368 187174 492688 187206
rect 492368 186938 492410 187174
rect 492646 186938 492688 187174
rect 492368 186854 492688 186938
rect 492368 186618 492410 186854
rect 492646 186618 492688 186854
rect 492368 186586 492688 186618
rect 523088 187174 523408 187206
rect 523088 186938 523130 187174
rect 523366 186938 523408 187174
rect 523088 186854 523408 186938
rect 523088 186618 523130 186854
rect 523366 186618 523408 186854
rect 523088 186586 523408 186618
rect 553808 187174 554128 187206
rect 553808 186938 553850 187174
rect 554086 186938 554128 187174
rect 553808 186854 554128 186938
rect 553808 186618 553850 186854
rect 554086 186618 554128 186854
rect 553808 186586 554128 186618
rect 16208 183454 16528 183486
rect 16208 183218 16250 183454
rect 16486 183218 16528 183454
rect 16208 183134 16528 183218
rect 16208 182898 16250 183134
rect 16486 182898 16528 183134
rect 16208 182866 16528 182898
rect 46928 183454 47248 183486
rect 46928 183218 46970 183454
rect 47206 183218 47248 183454
rect 46928 183134 47248 183218
rect 46928 182898 46970 183134
rect 47206 182898 47248 183134
rect 46928 182866 47248 182898
rect 77648 183454 77968 183486
rect 77648 183218 77690 183454
rect 77926 183218 77968 183454
rect 77648 183134 77968 183218
rect 77648 182898 77690 183134
rect 77926 182898 77968 183134
rect 77648 182866 77968 182898
rect 108368 183454 108688 183486
rect 108368 183218 108410 183454
rect 108646 183218 108688 183454
rect 108368 183134 108688 183218
rect 108368 182898 108410 183134
rect 108646 182898 108688 183134
rect 108368 182866 108688 182898
rect 139088 183454 139408 183486
rect 139088 183218 139130 183454
rect 139366 183218 139408 183454
rect 139088 183134 139408 183218
rect 139088 182898 139130 183134
rect 139366 182898 139408 183134
rect 139088 182866 139408 182898
rect 169808 183454 170128 183486
rect 169808 183218 169850 183454
rect 170086 183218 170128 183454
rect 169808 183134 170128 183218
rect 169808 182898 169850 183134
rect 170086 182898 170128 183134
rect 169808 182866 170128 182898
rect 200528 183454 200848 183486
rect 200528 183218 200570 183454
rect 200806 183218 200848 183454
rect 200528 183134 200848 183218
rect 200528 182898 200570 183134
rect 200806 182898 200848 183134
rect 200528 182866 200848 182898
rect 231248 183454 231568 183486
rect 231248 183218 231290 183454
rect 231526 183218 231568 183454
rect 231248 183134 231568 183218
rect 231248 182898 231290 183134
rect 231526 182898 231568 183134
rect 231248 182866 231568 182898
rect 261968 183454 262288 183486
rect 261968 183218 262010 183454
rect 262246 183218 262288 183454
rect 261968 183134 262288 183218
rect 261968 182898 262010 183134
rect 262246 182898 262288 183134
rect 261968 182866 262288 182898
rect 292688 183454 293008 183486
rect 292688 183218 292730 183454
rect 292966 183218 293008 183454
rect 292688 183134 293008 183218
rect 292688 182898 292730 183134
rect 292966 182898 293008 183134
rect 292688 182866 293008 182898
rect 323408 183454 323728 183486
rect 323408 183218 323450 183454
rect 323686 183218 323728 183454
rect 323408 183134 323728 183218
rect 323408 182898 323450 183134
rect 323686 182898 323728 183134
rect 323408 182866 323728 182898
rect 354128 183454 354448 183486
rect 354128 183218 354170 183454
rect 354406 183218 354448 183454
rect 354128 183134 354448 183218
rect 354128 182898 354170 183134
rect 354406 182898 354448 183134
rect 354128 182866 354448 182898
rect 384848 183454 385168 183486
rect 384848 183218 384890 183454
rect 385126 183218 385168 183454
rect 384848 183134 385168 183218
rect 384848 182898 384890 183134
rect 385126 182898 385168 183134
rect 384848 182866 385168 182898
rect 415568 183454 415888 183486
rect 415568 183218 415610 183454
rect 415846 183218 415888 183454
rect 415568 183134 415888 183218
rect 415568 182898 415610 183134
rect 415846 182898 415888 183134
rect 415568 182866 415888 182898
rect 446288 183454 446608 183486
rect 446288 183218 446330 183454
rect 446566 183218 446608 183454
rect 446288 183134 446608 183218
rect 446288 182898 446330 183134
rect 446566 182898 446608 183134
rect 446288 182866 446608 182898
rect 477008 183454 477328 183486
rect 477008 183218 477050 183454
rect 477286 183218 477328 183454
rect 477008 183134 477328 183218
rect 477008 182898 477050 183134
rect 477286 182898 477328 183134
rect 477008 182866 477328 182898
rect 507728 183454 508048 183486
rect 507728 183218 507770 183454
rect 508006 183218 508048 183454
rect 507728 183134 508048 183218
rect 507728 182898 507770 183134
rect 508006 182898 508048 183134
rect 507728 182866 508048 182898
rect 538448 183454 538768 183486
rect 538448 183218 538490 183454
rect 538726 183218 538768 183454
rect 538448 183134 538768 183218
rect 538448 182898 538490 183134
rect 538726 182898 538768 183134
rect 538448 182866 538768 182898
rect 9234 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 9854 154894
rect 9234 154574 9854 154658
rect 9234 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 9854 154574
rect 9234 118894 9854 154338
rect 567834 173494 568454 208938
rect 567834 173258 567866 173494
rect 568102 173258 568186 173494
rect 568422 173258 568454 173494
rect 567834 173174 568454 173258
rect 567834 172938 567866 173174
rect 568102 172938 568186 173174
rect 568422 172938 568454 173174
rect 31568 151174 31888 151206
rect 31568 150938 31610 151174
rect 31846 150938 31888 151174
rect 31568 150854 31888 150938
rect 31568 150618 31610 150854
rect 31846 150618 31888 150854
rect 31568 150586 31888 150618
rect 62288 151174 62608 151206
rect 62288 150938 62330 151174
rect 62566 150938 62608 151174
rect 62288 150854 62608 150938
rect 62288 150618 62330 150854
rect 62566 150618 62608 150854
rect 62288 150586 62608 150618
rect 93008 151174 93328 151206
rect 93008 150938 93050 151174
rect 93286 150938 93328 151174
rect 93008 150854 93328 150938
rect 93008 150618 93050 150854
rect 93286 150618 93328 150854
rect 93008 150586 93328 150618
rect 123728 151174 124048 151206
rect 123728 150938 123770 151174
rect 124006 150938 124048 151174
rect 123728 150854 124048 150938
rect 123728 150618 123770 150854
rect 124006 150618 124048 150854
rect 123728 150586 124048 150618
rect 154448 151174 154768 151206
rect 154448 150938 154490 151174
rect 154726 150938 154768 151174
rect 154448 150854 154768 150938
rect 154448 150618 154490 150854
rect 154726 150618 154768 150854
rect 154448 150586 154768 150618
rect 185168 151174 185488 151206
rect 185168 150938 185210 151174
rect 185446 150938 185488 151174
rect 185168 150854 185488 150938
rect 185168 150618 185210 150854
rect 185446 150618 185488 150854
rect 185168 150586 185488 150618
rect 215888 151174 216208 151206
rect 215888 150938 215930 151174
rect 216166 150938 216208 151174
rect 215888 150854 216208 150938
rect 215888 150618 215930 150854
rect 216166 150618 216208 150854
rect 215888 150586 216208 150618
rect 246608 151174 246928 151206
rect 246608 150938 246650 151174
rect 246886 150938 246928 151174
rect 246608 150854 246928 150938
rect 246608 150618 246650 150854
rect 246886 150618 246928 150854
rect 246608 150586 246928 150618
rect 277328 151174 277648 151206
rect 277328 150938 277370 151174
rect 277606 150938 277648 151174
rect 277328 150854 277648 150938
rect 277328 150618 277370 150854
rect 277606 150618 277648 150854
rect 277328 150586 277648 150618
rect 308048 151174 308368 151206
rect 308048 150938 308090 151174
rect 308326 150938 308368 151174
rect 308048 150854 308368 150938
rect 308048 150618 308090 150854
rect 308326 150618 308368 150854
rect 308048 150586 308368 150618
rect 338768 151174 339088 151206
rect 338768 150938 338810 151174
rect 339046 150938 339088 151174
rect 338768 150854 339088 150938
rect 338768 150618 338810 150854
rect 339046 150618 339088 150854
rect 338768 150586 339088 150618
rect 369488 151174 369808 151206
rect 369488 150938 369530 151174
rect 369766 150938 369808 151174
rect 369488 150854 369808 150938
rect 369488 150618 369530 150854
rect 369766 150618 369808 150854
rect 369488 150586 369808 150618
rect 400208 151174 400528 151206
rect 400208 150938 400250 151174
rect 400486 150938 400528 151174
rect 400208 150854 400528 150938
rect 400208 150618 400250 150854
rect 400486 150618 400528 150854
rect 400208 150586 400528 150618
rect 430928 151174 431248 151206
rect 430928 150938 430970 151174
rect 431206 150938 431248 151174
rect 430928 150854 431248 150938
rect 430928 150618 430970 150854
rect 431206 150618 431248 150854
rect 430928 150586 431248 150618
rect 461648 151174 461968 151206
rect 461648 150938 461690 151174
rect 461926 150938 461968 151174
rect 461648 150854 461968 150938
rect 461648 150618 461690 150854
rect 461926 150618 461968 150854
rect 461648 150586 461968 150618
rect 492368 151174 492688 151206
rect 492368 150938 492410 151174
rect 492646 150938 492688 151174
rect 492368 150854 492688 150938
rect 492368 150618 492410 150854
rect 492646 150618 492688 150854
rect 492368 150586 492688 150618
rect 523088 151174 523408 151206
rect 523088 150938 523130 151174
rect 523366 150938 523408 151174
rect 523088 150854 523408 150938
rect 523088 150618 523130 150854
rect 523366 150618 523408 150854
rect 523088 150586 523408 150618
rect 553808 151174 554128 151206
rect 553808 150938 553850 151174
rect 554086 150938 554128 151174
rect 553808 150854 554128 150938
rect 553808 150618 553850 150854
rect 554086 150618 554128 150854
rect 553808 150586 554128 150618
rect 16208 147454 16528 147486
rect 16208 147218 16250 147454
rect 16486 147218 16528 147454
rect 16208 147134 16528 147218
rect 16208 146898 16250 147134
rect 16486 146898 16528 147134
rect 16208 146866 16528 146898
rect 46928 147454 47248 147486
rect 46928 147218 46970 147454
rect 47206 147218 47248 147454
rect 46928 147134 47248 147218
rect 46928 146898 46970 147134
rect 47206 146898 47248 147134
rect 46928 146866 47248 146898
rect 77648 147454 77968 147486
rect 77648 147218 77690 147454
rect 77926 147218 77968 147454
rect 77648 147134 77968 147218
rect 77648 146898 77690 147134
rect 77926 146898 77968 147134
rect 77648 146866 77968 146898
rect 108368 147454 108688 147486
rect 108368 147218 108410 147454
rect 108646 147218 108688 147454
rect 108368 147134 108688 147218
rect 108368 146898 108410 147134
rect 108646 146898 108688 147134
rect 108368 146866 108688 146898
rect 139088 147454 139408 147486
rect 139088 147218 139130 147454
rect 139366 147218 139408 147454
rect 139088 147134 139408 147218
rect 139088 146898 139130 147134
rect 139366 146898 139408 147134
rect 139088 146866 139408 146898
rect 169808 147454 170128 147486
rect 169808 147218 169850 147454
rect 170086 147218 170128 147454
rect 169808 147134 170128 147218
rect 169808 146898 169850 147134
rect 170086 146898 170128 147134
rect 169808 146866 170128 146898
rect 200528 147454 200848 147486
rect 200528 147218 200570 147454
rect 200806 147218 200848 147454
rect 200528 147134 200848 147218
rect 200528 146898 200570 147134
rect 200806 146898 200848 147134
rect 200528 146866 200848 146898
rect 231248 147454 231568 147486
rect 231248 147218 231290 147454
rect 231526 147218 231568 147454
rect 231248 147134 231568 147218
rect 231248 146898 231290 147134
rect 231526 146898 231568 147134
rect 231248 146866 231568 146898
rect 261968 147454 262288 147486
rect 261968 147218 262010 147454
rect 262246 147218 262288 147454
rect 261968 147134 262288 147218
rect 261968 146898 262010 147134
rect 262246 146898 262288 147134
rect 261968 146866 262288 146898
rect 292688 147454 293008 147486
rect 292688 147218 292730 147454
rect 292966 147218 293008 147454
rect 292688 147134 293008 147218
rect 292688 146898 292730 147134
rect 292966 146898 293008 147134
rect 292688 146866 293008 146898
rect 323408 147454 323728 147486
rect 323408 147218 323450 147454
rect 323686 147218 323728 147454
rect 323408 147134 323728 147218
rect 323408 146898 323450 147134
rect 323686 146898 323728 147134
rect 323408 146866 323728 146898
rect 354128 147454 354448 147486
rect 354128 147218 354170 147454
rect 354406 147218 354448 147454
rect 354128 147134 354448 147218
rect 354128 146898 354170 147134
rect 354406 146898 354448 147134
rect 354128 146866 354448 146898
rect 384848 147454 385168 147486
rect 384848 147218 384890 147454
rect 385126 147218 385168 147454
rect 384848 147134 385168 147218
rect 384848 146898 384890 147134
rect 385126 146898 385168 147134
rect 384848 146866 385168 146898
rect 415568 147454 415888 147486
rect 415568 147218 415610 147454
rect 415846 147218 415888 147454
rect 415568 147134 415888 147218
rect 415568 146898 415610 147134
rect 415846 146898 415888 147134
rect 415568 146866 415888 146898
rect 446288 147454 446608 147486
rect 446288 147218 446330 147454
rect 446566 147218 446608 147454
rect 446288 147134 446608 147218
rect 446288 146898 446330 147134
rect 446566 146898 446608 147134
rect 446288 146866 446608 146898
rect 477008 147454 477328 147486
rect 477008 147218 477050 147454
rect 477286 147218 477328 147454
rect 477008 147134 477328 147218
rect 477008 146898 477050 147134
rect 477286 146898 477328 147134
rect 477008 146866 477328 146898
rect 507728 147454 508048 147486
rect 507728 147218 507770 147454
rect 508006 147218 508048 147454
rect 507728 147134 508048 147218
rect 507728 146898 507770 147134
rect 508006 146898 508048 147134
rect 507728 146866 508048 146898
rect 538448 147454 538768 147486
rect 538448 147218 538490 147454
rect 538726 147218 538768 147454
rect 538448 147134 538768 147218
rect 538448 146898 538490 147134
rect 538726 146898 538768 147134
rect 538448 146866 538768 146898
rect 9234 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 9854 118894
rect 9234 118574 9854 118658
rect 9234 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 9854 118574
rect 9234 82894 9854 118338
rect 567834 137494 568454 172938
rect 567834 137258 567866 137494
rect 568102 137258 568186 137494
rect 568422 137258 568454 137494
rect 567834 137174 568454 137258
rect 567834 136938 567866 137174
rect 568102 136938 568186 137174
rect 568422 136938 568454 137174
rect 31568 115174 31888 115206
rect 31568 114938 31610 115174
rect 31846 114938 31888 115174
rect 31568 114854 31888 114938
rect 31568 114618 31610 114854
rect 31846 114618 31888 114854
rect 31568 114586 31888 114618
rect 62288 115174 62608 115206
rect 62288 114938 62330 115174
rect 62566 114938 62608 115174
rect 62288 114854 62608 114938
rect 62288 114618 62330 114854
rect 62566 114618 62608 114854
rect 62288 114586 62608 114618
rect 93008 115174 93328 115206
rect 93008 114938 93050 115174
rect 93286 114938 93328 115174
rect 93008 114854 93328 114938
rect 93008 114618 93050 114854
rect 93286 114618 93328 114854
rect 93008 114586 93328 114618
rect 123728 115174 124048 115206
rect 123728 114938 123770 115174
rect 124006 114938 124048 115174
rect 123728 114854 124048 114938
rect 123728 114618 123770 114854
rect 124006 114618 124048 114854
rect 123728 114586 124048 114618
rect 154448 115174 154768 115206
rect 154448 114938 154490 115174
rect 154726 114938 154768 115174
rect 154448 114854 154768 114938
rect 154448 114618 154490 114854
rect 154726 114618 154768 114854
rect 154448 114586 154768 114618
rect 185168 115174 185488 115206
rect 185168 114938 185210 115174
rect 185446 114938 185488 115174
rect 185168 114854 185488 114938
rect 185168 114618 185210 114854
rect 185446 114618 185488 114854
rect 185168 114586 185488 114618
rect 215888 115174 216208 115206
rect 215888 114938 215930 115174
rect 216166 114938 216208 115174
rect 215888 114854 216208 114938
rect 215888 114618 215930 114854
rect 216166 114618 216208 114854
rect 215888 114586 216208 114618
rect 246608 115174 246928 115206
rect 246608 114938 246650 115174
rect 246886 114938 246928 115174
rect 246608 114854 246928 114938
rect 246608 114618 246650 114854
rect 246886 114618 246928 114854
rect 246608 114586 246928 114618
rect 277328 115174 277648 115206
rect 277328 114938 277370 115174
rect 277606 114938 277648 115174
rect 277328 114854 277648 114938
rect 277328 114618 277370 114854
rect 277606 114618 277648 114854
rect 277328 114586 277648 114618
rect 308048 115174 308368 115206
rect 308048 114938 308090 115174
rect 308326 114938 308368 115174
rect 308048 114854 308368 114938
rect 308048 114618 308090 114854
rect 308326 114618 308368 114854
rect 308048 114586 308368 114618
rect 338768 115174 339088 115206
rect 338768 114938 338810 115174
rect 339046 114938 339088 115174
rect 338768 114854 339088 114938
rect 338768 114618 338810 114854
rect 339046 114618 339088 114854
rect 338768 114586 339088 114618
rect 369488 115174 369808 115206
rect 369488 114938 369530 115174
rect 369766 114938 369808 115174
rect 369488 114854 369808 114938
rect 369488 114618 369530 114854
rect 369766 114618 369808 114854
rect 369488 114586 369808 114618
rect 400208 115174 400528 115206
rect 400208 114938 400250 115174
rect 400486 114938 400528 115174
rect 400208 114854 400528 114938
rect 400208 114618 400250 114854
rect 400486 114618 400528 114854
rect 400208 114586 400528 114618
rect 430928 115174 431248 115206
rect 430928 114938 430970 115174
rect 431206 114938 431248 115174
rect 430928 114854 431248 114938
rect 430928 114618 430970 114854
rect 431206 114618 431248 114854
rect 430928 114586 431248 114618
rect 461648 115174 461968 115206
rect 461648 114938 461690 115174
rect 461926 114938 461968 115174
rect 461648 114854 461968 114938
rect 461648 114618 461690 114854
rect 461926 114618 461968 114854
rect 461648 114586 461968 114618
rect 492368 115174 492688 115206
rect 492368 114938 492410 115174
rect 492646 114938 492688 115174
rect 492368 114854 492688 114938
rect 492368 114618 492410 114854
rect 492646 114618 492688 114854
rect 492368 114586 492688 114618
rect 523088 115174 523408 115206
rect 523088 114938 523130 115174
rect 523366 114938 523408 115174
rect 523088 114854 523408 114938
rect 523088 114618 523130 114854
rect 523366 114618 523408 114854
rect 523088 114586 523408 114618
rect 553808 115174 554128 115206
rect 553808 114938 553850 115174
rect 554086 114938 554128 115174
rect 553808 114854 554128 114938
rect 553808 114618 553850 114854
rect 554086 114618 554128 114854
rect 553808 114586 554128 114618
rect 16208 111454 16528 111486
rect 16208 111218 16250 111454
rect 16486 111218 16528 111454
rect 16208 111134 16528 111218
rect 16208 110898 16250 111134
rect 16486 110898 16528 111134
rect 16208 110866 16528 110898
rect 46928 111454 47248 111486
rect 46928 111218 46970 111454
rect 47206 111218 47248 111454
rect 46928 111134 47248 111218
rect 46928 110898 46970 111134
rect 47206 110898 47248 111134
rect 46928 110866 47248 110898
rect 77648 111454 77968 111486
rect 77648 111218 77690 111454
rect 77926 111218 77968 111454
rect 77648 111134 77968 111218
rect 77648 110898 77690 111134
rect 77926 110898 77968 111134
rect 77648 110866 77968 110898
rect 108368 111454 108688 111486
rect 108368 111218 108410 111454
rect 108646 111218 108688 111454
rect 108368 111134 108688 111218
rect 108368 110898 108410 111134
rect 108646 110898 108688 111134
rect 108368 110866 108688 110898
rect 139088 111454 139408 111486
rect 139088 111218 139130 111454
rect 139366 111218 139408 111454
rect 139088 111134 139408 111218
rect 139088 110898 139130 111134
rect 139366 110898 139408 111134
rect 139088 110866 139408 110898
rect 169808 111454 170128 111486
rect 169808 111218 169850 111454
rect 170086 111218 170128 111454
rect 169808 111134 170128 111218
rect 169808 110898 169850 111134
rect 170086 110898 170128 111134
rect 169808 110866 170128 110898
rect 200528 111454 200848 111486
rect 200528 111218 200570 111454
rect 200806 111218 200848 111454
rect 200528 111134 200848 111218
rect 200528 110898 200570 111134
rect 200806 110898 200848 111134
rect 200528 110866 200848 110898
rect 231248 111454 231568 111486
rect 231248 111218 231290 111454
rect 231526 111218 231568 111454
rect 231248 111134 231568 111218
rect 231248 110898 231290 111134
rect 231526 110898 231568 111134
rect 231248 110866 231568 110898
rect 261968 111454 262288 111486
rect 261968 111218 262010 111454
rect 262246 111218 262288 111454
rect 261968 111134 262288 111218
rect 261968 110898 262010 111134
rect 262246 110898 262288 111134
rect 261968 110866 262288 110898
rect 292688 111454 293008 111486
rect 292688 111218 292730 111454
rect 292966 111218 293008 111454
rect 292688 111134 293008 111218
rect 292688 110898 292730 111134
rect 292966 110898 293008 111134
rect 292688 110866 293008 110898
rect 323408 111454 323728 111486
rect 323408 111218 323450 111454
rect 323686 111218 323728 111454
rect 323408 111134 323728 111218
rect 323408 110898 323450 111134
rect 323686 110898 323728 111134
rect 323408 110866 323728 110898
rect 354128 111454 354448 111486
rect 354128 111218 354170 111454
rect 354406 111218 354448 111454
rect 354128 111134 354448 111218
rect 354128 110898 354170 111134
rect 354406 110898 354448 111134
rect 354128 110866 354448 110898
rect 384848 111454 385168 111486
rect 384848 111218 384890 111454
rect 385126 111218 385168 111454
rect 384848 111134 385168 111218
rect 384848 110898 384890 111134
rect 385126 110898 385168 111134
rect 384848 110866 385168 110898
rect 415568 111454 415888 111486
rect 415568 111218 415610 111454
rect 415846 111218 415888 111454
rect 415568 111134 415888 111218
rect 415568 110898 415610 111134
rect 415846 110898 415888 111134
rect 415568 110866 415888 110898
rect 446288 111454 446608 111486
rect 446288 111218 446330 111454
rect 446566 111218 446608 111454
rect 446288 111134 446608 111218
rect 446288 110898 446330 111134
rect 446566 110898 446608 111134
rect 446288 110866 446608 110898
rect 477008 111454 477328 111486
rect 477008 111218 477050 111454
rect 477286 111218 477328 111454
rect 477008 111134 477328 111218
rect 477008 110898 477050 111134
rect 477286 110898 477328 111134
rect 477008 110866 477328 110898
rect 507728 111454 508048 111486
rect 507728 111218 507770 111454
rect 508006 111218 508048 111454
rect 507728 111134 508048 111218
rect 507728 110898 507770 111134
rect 508006 110898 508048 111134
rect 507728 110866 508048 110898
rect 538448 111454 538768 111486
rect 538448 111218 538490 111454
rect 538726 111218 538768 111454
rect 538448 111134 538768 111218
rect 538448 110898 538490 111134
rect 538726 110898 538768 111134
rect 538448 110866 538768 110898
rect 9234 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 9854 82894
rect 9234 82574 9854 82658
rect 9234 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 9854 82574
rect 9234 46894 9854 82338
rect 567834 101494 568454 136938
rect 567834 101258 567866 101494
rect 568102 101258 568186 101494
rect 568422 101258 568454 101494
rect 567834 101174 568454 101258
rect 567834 100938 567866 101174
rect 568102 100938 568186 101174
rect 568422 100938 568454 101174
rect 31568 79174 31888 79206
rect 31568 78938 31610 79174
rect 31846 78938 31888 79174
rect 31568 78854 31888 78938
rect 31568 78618 31610 78854
rect 31846 78618 31888 78854
rect 31568 78586 31888 78618
rect 62288 79174 62608 79206
rect 62288 78938 62330 79174
rect 62566 78938 62608 79174
rect 62288 78854 62608 78938
rect 62288 78618 62330 78854
rect 62566 78618 62608 78854
rect 62288 78586 62608 78618
rect 93008 79174 93328 79206
rect 93008 78938 93050 79174
rect 93286 78938 93328 79174
rect 93008 78854 93328 78938
rect 93008 78618 93050 78854
rect 93286 78618 93328 78854
rect 93008 78586 93328 78618
rect 123728 79174 124048 79206
rect 123728 78938 123770 79174
rect 124006 78938 124048 79174
rect 123728 78854 124048 78938
rect 123728 78618 123770 78854
rect 124006 78618 124048 78854
rect 123728 78586 124048 78618
rect 154448 79174 154768 79206
rect 154448 78938 154490 79174
rect 154726 78938 154768 79174
rect 154448 78854 154768 78938
rect 154448 78618 154490 78854
rect 154726 78618 154768 78854
rect 154448 78586 154768 78618
rect 185168 79174 185488 79206
rect 185168 78938 185210 79174
rect 185446 78938 185488 79174
rect 185168 78854 185488 78938
rect 185168 78618 185210 78854
rect 185446 78618 185488 78854
rect 185168 78586 185488 78618
rect 215888 79174 216208 79206
rect 215888 78938 215930 79174
rect 216166 78938 216208 79174
rect 215888 78854 216208 78938
rect 215888 78618 215930 78854
rect 216166 78618 216208 78854
rect 215888 78586 216208 78618
rect 246608 79174 246928 79206
rect 246608 78938 246650 79174
rect 246886 78938 246928 79174
rect 246608 78854 246928 78938
rect 246608 78618 246650 78854
rect 246886 78618 246928 78854
rect 246608 78586 246928 78618
rect 277328 79174 277648 79206
rect 277328 78938 277370 79174
rect 277606 78938 277648 79174
rect 277328 78854 277648 78938
rect 277328 78618 277370 78854
rect 277606 78618 277648 78854
rect 277328 78586 277648 78618
rect 308048 79174 308368 79206
rect 308048 78938 308090 79174
rect 308326 78938 308368 79174
rect 308048 78854 308368 78938
rect 308048 78618 308090 78854
rect 308326 78618 308368 78854
rect 308048 78586 308368 78618
rect 338768 79174 339088 79206
rect 338768 78938 338810 79174
rect 339046 78938 339088 79174
rect 338768 78854 339088 78938
rect 338768 78618 338810 78854
rect 339046 78618 339088 78854
rect 338768 78586 339088 78618
rect 369488 79174 369808 79206
rect 369488 78938 369530 79174
rect 369766 78938 369808 79174
rect 369488 78854 369808 78938
rect 369488 78618 369530 78854
rect 369766 78618 369808 78854
rect 369488 78586 369808 78618
rect 400208 79174 400528 79206
rect 400208 78938 400250 79174
rect 400486 78938 400528 79174
rect 400208 78854 400528 78938
rect 400208 78618 400250 78854
rect 400486 78618 400528 78854
rect 400208 78586 400528 78618
rect 430928 79174 431248 79206
rect 430928 78938 430970 79174
rect 431206 78938 431248 79174
rect 430928 78854 431248 78938
rect 430928 78618 430970 78854
rect 431206 78618 431248 78854
rect 430928 78586 431248 78618
rect 461648 79174 461968 79206
rect 461648 78938 461690 79174
rect 461926 78938 461968 79174
rect 461648 78854 461968 78938
rect 461648 78618 461690 78854
rect 461926 78618 461968 78854
rect 461648 78586 461968 78618
rect 492368 79174 492688 79206
rect 492368 78938 492410 79174
rect 492646 78938 492688 79174
rect 492368 78854 492688 78938
rect 492368 78618 492410 78854
rect 492646 78618 492688 78854
rect 492368 78586 492688 78618
rect 523088 79174 523408 79206
rect 523088 78938 523130 79174
rect 523366 78938 523408 79174
rect 523088 78854 523408 78938
rect 523088 78618 523130 78854
rect 523366 78618 523408 78854
rect 523088 78586 523408 78618
rect 553808 79174 554128 79206
rect 553808 78938 553850 79174
rect 554086 78938 554128 79174
rect 553808 78854 554128 78938
rect 553808 78618 553850 78854
rect 554086 78618 554128 78854
rect 553808 78586 554128 78618
rect 16208 75454 16528 75486
rect 16208 75218 16250 75454
rect 16486 75218 16528 75454
rect 16208 75134 16528 75218
rect 16208 74898 16250 75134
rect 16486 74898 16528 75134
rect 16208 74866 16528 74898
rect 46928 75454 47248 75486
rect 46928 75218 46970 75454
rect 47206 75218 47248 75454
rect 46928 75134 47248 75218
rect 46928 74898 46970 75134
rect 47206 74898 47248 75134
rect 46928 74866 47248 74898
rect 77648 75454 77968 75486
rect 77648 75218 77690 75454
rect 77926 75218 77968 75454
rect 77648 75134 77968 75218
rect 77648 74898 77690 75134
rect 77926 74898 77968 75134
rect 77648 74866 77968 74898
rect 108368 75454 108688 75486
rect 108368 75218 108410 75454
rect 108646 75218 108688 75454
rect 108368 75134 108688 75218
rect 108368 74898 108410 75134
rect 108646 74898 108688 75134
rect 108368 74866 108688 74898
rect 139088 75454 139408 75486
rect 139088 75218 139130 75454
rect 139366 75218 139408 75454
rect 139088 75134 139408 75218
rect 139088 74898 139130 75134
rect 139366 74898 139408 75134
rect 139088 74866 139408 74898
rect 169808 75454 170128 75486
rect 169808 75218 169850 75454
rect 170086 75218 170128 75454
rect 169808 75134 170128 75218
rect 169808 74898 169850 75134
rect 170086 74898 170128 75134
rect 169808 74866 170128 74898
rect 200528 75454 200848 75486
rect 200528 75218 200570 75454
rect 200806 75218 200848 75454
rect 200528 75134 200848 75218
rect 200528 74898 200570 75134
rect 200806 74898 200848 75134
rect 200528 74866 200848 74898
rect 231248 75454 231568 75486
rect 231248 75218 231290 75454
rect 231526 75218 231568 75454
rect 231248 75134 231568 75218
rect 231248 74898 231290 75134
rect 231526 74898 231568 75134
rect 231248 74866 231568 74898
rect 261968 75454 262288 75486
rect 261968 75218 262010 75454
rect 262246 75218 262288 75454
rect 261968 75134 262288 75218
rect 261968 74898 262010 75134
rect 262246 74898 262288 75134
rect 261968 74866 262288 74898
rect 292688 75454 293008 75486
rect 292688 75218 292730 75454
rect 292966 75218 293008 75454
rect 292688 75134 293008 75218
rect 292688 74898 292730 75134
rect 292966 74898 293008 75134
rect 292688 74866 293008 74898
rect 323408 75454 323728 75486
rect 323408 75218 323450 75454
rect 323686 75218 323728 75454
rect 323408 75134 323728 75218
rect 323408 74898 323450 75134
rect 323686 74898 323728 75134
rect 323408 74866 323728 74898
rect 354128 75454 354448 75486
rect 354128 75218 354170 75454
rect 354406 75218 354448 75454
rect 354128 75134 354448 75218
rect 354128 74898 354170 75134
rect 354406 74898 354448 75134
rect 354128 74866 354448 74898
rect 384848 75454 385168 75486
rect 384848 75218 384890 75454
rect 385126 75218 385168 75454
rect 384848 75134 385168 75218
rect 384848 74898 384890 75134
rect 385126 74898 385168 75134
rect 384848 74866 385168 74898
rect 415568 75454 415888 75486
rect 415568 75218 415610 75454
rect 415846 75218 415888 75454
rect 415568 75134 415888 75218
rect 415568 74898 415610 75134
rect 415846 74898 415888 75134
rect 415568 74866 415888 74898
rect 446288 75454 446608 75486
rect 446288 75218 446330 75454
rect 446566 75218 446608 75454
rect 446288 75134 446608 75218
rect 446288 74898 446330 75134
rect 446566 74898 446608 75134
rect 446288 74866 446608 74898
rect 477008 75454 477328 75486
rect 477008 75218 477050 75454
rect 477286 75218 477328 75454
rect 477008 75134 477328 75218
rect 477008 74898 477050 75134
rect 477286 74898 477328 75134
rect 477008 74866 477328 74898
rect 507728 75454 508048 75486
rect 507728 75218 507770 75454
rect 508006 75218 508048 75454
rect 507728 75134 508048 75218
rect 507728 74898 507770 75134
rect 508006 74898 508048 75134
rect 507728 74866 508048 74898
rect 538448 75454 538768 75486
rect 538448 75218 538490 75454
rect 538726 75218 538768 75454
rect 538448 75134 538768 75218
rect 538448 74898 538490 75134
rect 538726 74898 538768 75134
rect 538448 74866 538768 74898
rect 9234 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 9854 46894
rect 9234 46574 9854 46658
rect 9234 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 9854 46574
rect 9234 10894 9854 46338
rect 567834 65494 568454 100938
rect 567834 65258 567866 65494
rect 568102 65258 568186 65494
rect 568422 65258 568454 65494
rect 567834 65174 568454 65258
rect 567834 64938 567866 65174
rect 568102 64938 568186 65174
rect 568422 64938 568454 65174
rect 31568 43174 31888 43206
rect 31568 42938 31610 43174
rect 31846 42938 31888 43174
rect 31568 42854 31888 42938
rect 31568 42618 31610 42854
rect 31846 42618 31888 42854
rect 31568 42586 31888 42618
rect 62288 43174 62608 43206
rect 62288 42938 62330 43174
rect 62566 42938 62608 43174
rect 62288 42854 62608 42938
rect 62288 42618 62330 42854
rect 62566 42618 62608 42854
rect 62288 42586 62608 42618
rect 93008 43174 93328 43206
rect 93008 42938 93050 43174
rect 93286 42938 93328 43174
rect 93008 42854 93328 42938
rect 93008 42618 93050 42854
rect 93286 42618 93328 42854
rect 93008 42586 93328 42618
rect 123728 43174 124048 43206
rect 123728 42938 123770 43174
rect 124006 42938 124048 43174
rect 123728 42854 124048 42938
rect 123728 42618 123770 42854
rect 124006 42618 124048 42854
rect 123728 42586 124048 42618
rect 154448 43174 154768 43206
rect 154448 42938 154490 43174
rect 154726 42938 154768 43174
rect 154448 42854 154768 42938
rect 154448 42618 154490 42854
rect 154726 42618 154768 42854
rect 154448 42586 154768 42618
rect 185168 43174 185488 43206
rect 185168 42938 185210 43174
rect 185446 42938 185488 43174
rect 185168 42854 185488 42938
rect 185168 42618 185210 42854
rect 185446 42618 185488 42854
rect 185168 42586 185488 42618
rect 215888 43174 216208 43206
rect 215888 42938 215930 43174
rect 216166 42938 216208 43174
rect 215888 42854 216208 42938
rect 215888 42618 215930 42854
rect 216166 42618 216208 42854
rect 215888 42586 216208 42618
rect 246608 43174 246928 43206
rect 246608 42938 246650 43174
rect 246886 42938 246928 43174
rect 246608 42854 246928 42938
rect 246608 42618 246650 42854
rect 246886 42618 246928 42854
rect 246608 42586 246928 42618
rect 277328 43174 277648 43206
rect 277328 42938 277370 43174
rect 277606 42938 277648 43174
rect 277328 42854 277648 42938
rect 277328 42618 277370 42854
rect 277606 42618 277648 42854
rect 277328 42586 277648 42618
rect 308048 43174 308368 43206
rect 308048 42938 308090 43174
rect 308326 42938 308368 43174
rect 308048 42854 308368 42938
rect 308048 42618 308090 42854
rect 308326 42618 308368 42854
rect 308048 42586 308368 42618
rect 338768 43174 339088 43206
rect 338768 42938 338810 43174
rect 339046 42938 339088 43174
rect 338768 42854 339088 42938
rect 338768 42618 338810 42854
rect 339046 42618 339088 42854
rect 338768 42586 339088 42618
rect 369488 43174 369808 43206
rect 369488 42938 369530 43174
rect 369766 42938 369808 43174
rect 369488 42854 369808 42938
rect 369488 42618 369530 42854
rect 369766 42618 369808 42854
rect 369488 42586 369808 42618
rect 400208 43174 400528 43206
rect 400208 42938 400250 43174
rect 400486 42938 400528 43174
rect 400208 42854 400528 42938
rect 400208 42618 400250 42854
rect 400486 42618 400528 42854
rect 400208 42586 400528 42618
rect 430928 43174 431248 43206
rect 430928 42938 430970 43174
rect 431206 42938 431248 43174
rect 430928 42854 431248 42938
rect 430928 42618 430970 42854
rect 431206 42618 431248 42854
rect 430928 42586 431248 42618
rect 461648 43174 461968 43206
rect 461648 42938 461690 43174
rect 461926 42938 461968 43174
rect 461648 42854 461968 42938
rect 461648 42618 461690 42854
rect 461926 42618 461968 42854
rect 461648 42586 461968 42618
rect 492368 43174 492688 43206
rect 492368 42938 492410 43174
rect 492646 42938 492688 43174
rect 492368 42854 492688 42938
rect 492368 42618 492410 42854
rect 492646 42618 492688 42854
rect 492368 42586 492688 42618
rect 523088 43174 523408 43206
rect 523088 42938 523130 43174
rect 523366 42938 523408 43174
rect 523088 42854 523408 42938
rect 523088 42618 523130 42854
rect 523366 42618 523408 42854
rect 523088 42586 523408 42618
rect 553808 43174 554128 43206
rect 553808 42938 553850 43174
rect 554086 42938 554128 43174
rect 553808 42854 554128 42938
rect 553808 42618 553850 42854
rect 554086 42618 554128 42854
rect 553808 42586 554128 42618
rect 16208 39454 16528 39486
rect 16208 39218 16250 39454
rect 16486 39218 16528 39454
rect 16208 39134 16528 39218
rect 16208 38898 16250 39134
rect 16486 38898 16528 39134
rect 16208 38866 16528 38898
rect 46928 39454 47248 39486
rect 46928 39218 46970 39454
rect 47206 39218 47248 39454
rect 46928 39134 47248 39218
rect 46928 38898 46970 39134
rect 47206 38898 47248 39134
rect 46928 38866 47248 38898
rect 77648 39454 77968 39486
rect 77648 39218 77690 39454
rect 77926 39218 77968 39454
rect 77648 39134 77968 39218
rect 77648 38898 77690 39134
rect 77926 38898 77968 39134
rect 77648 38866 77968 38898
rect 108368 39454 108688 39486
rect 108368 39218 108410 39454
rect 108646 39218 108688 39454
rect 108368 39134 108688 39218
rect 108368 38898 108410 39134
rect 108646 38898 108688 39134
rect 108368 38866 108688 38898
rect 139088 39454 139408 39486
rect 139088 39218 139130 39454
rect 139366 39218 139408 39454
rect 139088 39134 139408 39218
rect 139088 38898 139130 39134
rect 139366 38898 139408 39134
rect 139088 38866 139408 38898
rect 169808 39454 170128 39486
rect 169808 39218 169850 39454
rect 170086 39218 170128 39454
rect 169808 39134 170128 39218
rect 169808 38898 169850 39134
rect 170086 38898 170128 39134
rect 169808 38866 170128 38898
rect 200528 39454 200848 39486
rect 200528 39218 200570 39454
rect 200806 39218 200848 39454
rect 200528 39134 200848 39218
rect 200528 38898 200570 39134
rect 200806 38898 200848 39134
rect 200528 38866 200848 38898
rect 231248 39454 231568 39486
rect 231248 39218 231290 39454
rect 231526 39218 231568 39454
rect 231248 39134 231568 39218
rect 231248 38898 231290 39134
rect 231526 38898 231568 39134
rect 231248 38866 231568 38898
rect 261968 39454 262288 39486
rect 261968 39218 262010 39454
rect 262246 39218 262288 39454
rect 261968 39134 262288 39218
rect 261968 38898 262010 39134
rect 262246 38898 262288 39134
rect 261968 38866 262288 38898
rect 292688 39454 293008 39486
rect 292688 39218 292730 39454
rect 292966 39218 293008 39454
rect 292688 39134 293008 39218
rect 292688 38898 292730 39134
rect 292966 38898 293008 39134
rect 292688 38866 293008 38898
rect 323408 39454 323728 39486
rect 323408 39218 323450 39454
rect 323686 39218 323728 39454
rect 323408 39134 323728 39218
rect 323408 38898 323450 39134
rect 323686 38898 323728 39134
rect 323408 38866 323728 38898
rect 354128 39454 354448 39486
rect 354128 39218 354170 39454
rect 354406 39218 354448 39454
rect 354128 39134 354448 39218
rect 354128 38898 354170 39134
rect 354406 38898 354448 39134
rect 354128 38866 354448 38898
rect 384848 39454 385168 39486
rect 384848 39218 384890 39454
rect 385126 39218 385168 39454
rect 384848 39134 385168 39218
rect 384848 38898 384890 39134
rect 385126 38898 385168 39134
rect 384848 38866 385168 38898
rect 415568 39454 415888 39486
rect 415568 39218 415610 39454
rect 415846 39218 415888 39454
rect 415568 39134 415888 39218
rect 415568 38898 415610 39134
rect 415846 38898 415888 39134
rect 415568 38866 415888 38898
rect 446288 39454 446608 39486
rect 446288 39218 446330 39454
rect 446566 39218 446608 39454
rect 446288 39134 446608 39218
rect 446288 38898 446330 39134
rect 446566 38898 446608 39134
rect 446288 38866 446608 38898
rect 477008 39454 477328 39486
rect 477008 39218 477050 39454
rect 477286 39218 477328 39454
rect 477008 39134 477328 39218
rect 477008 38898 477050 39134
rect 477286 38898 477328 39134
rect 477008 38866 477328 38898
rect 507728 39454 508048 39486
rect 507728 39218 507770 39454
rect 508006 39218 508048 39454
rect 507728 39134 508048 39218
rect 507728 38898 507770 39134
rect 508006 38898 508048 39134
rect 507728 38866 508048 38898
rect 538448 39454 538768 39486
rect 538448 39218 538490 39454
rect 538726 39218 538768 39454
rect 538448 39134 538768 39218
rect 538448 38898 538490 39134
rect 538726 38898 538768 39134
rect 538448 38866 538768 38898
rect 567834 29494 568454 64938
rect 567834 29258 567866 29494
rect 568102 29258 568186 29494
rect 568422 29258 568454 29494
rect 567834 29174 568454 29258
rect 567834 28938 567866 29174
rect 568102 28938 568186 29174
rect 568422 28938 568454 29174
rect 9234 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 9854 10894
rect 9234 10574 9854 10658
rect 9234 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 9854 10574
rect 9234 -2266 9854 10338
rect 9234 -2502 9266 -2266
rect 9502 -2502 9586 -2266
rect 9822 -2502 9854 -2266
rect 9234 -2586 9854 -2502
rect 9234 -2822 9266 -2586
rect 9502 -2822 9586 -2586
rect 9822 -2822 9854 -2586
rect 9234 -7654 9854 -2822
rect 37794 3454 38414 12559
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -7654 38414 -902
rect 41514 7174 42134 12559
rect 41514 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 42134 7174
rect 41514 6854 42134 6938
rect 41514 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 42134 6854
rect 41514 -1306 42134 6618
rect 41514 -1542 41546 -1306
rect 41782 -1542 41866 -1306
rect 42102 -1542 42134 -1306
rect 41514 -1626 42134 -1542
rect 41514 -1862 41546 -1626
rect 41782 -1862 41866 -1626
rect 42102 -1862 42134 -1626
rect 41514 -7654 42134 -1862
rect 45234 10894 45854 12559
rect 45234 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 45854 10894
rect 45234 10574 45854 10658
rect 45234 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 45854 10574
rect 45234 -2266 45854 10338
rect 45234 -2502 45266 -2266
rect 45502 -2502 45586 -2266
rect 45822 -2502 45854 -2266
rect 45234 -2586 45854 -2502
rect 45234 -2822 45266 -2586
rect 45502 -2822 45586 -2586
rect 45822 -2822 45854 -2586
rect 45234 -7654 45854 -2822
rect 73794 3454 74414 12559
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -7654 74414 -902
rect 77514 7174 78134 12068
rect 77514 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 78134 7174
rect 77514 6854 78134 6938
rect 77514 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 78134 6854
rect 77514 -1306 78134 6618
rect 77514 -1542 77546 -1306
rect 77782 -1542 77866 -1306
rect 78102 -1542 78134 -1306
rect 77514 -1626 78134 -1542
rect 77514 -1862 77546 -1626
rect 77782 -1862 77866 -1626
rect 78102 -1862 78134 -1626
rect 77514 -7654 78134 -1862
rect 81234 10894 81854 12559
rect 81234 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 81854 10894
rect 81234 10574 81854 10658
rect 81234 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 81854 10574
rect 81234 -2266 81854 10338
rect 81234 -2502 81266 -2266
rect 81502 -2502 81586 -2266
rect 81822 -2502 81854 -2266
rect 81234 -2586 81854 -2502
rect 81234 -2822 81266 -2586
rect 81502 -2822 81586 -2586
rect 81822 -2822 81854 -2586
rect 81234 -7654 81854 -2822
rect 109794 3454 110414 12559
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -7654 110414 -902
rect 113514 7174 114134 12559
rect 113514 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 114134 7174
rect 113514 6854 114134 6938
rect 113514 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 114134 6854
rect 113514 -1306 114134 6618
rect 113514 -1542 113546 -1306
rect 113782 -1542 113866 -1306
rect 114102 -1542 114134 -1306
rect 113514 -1626 114134 -1542
rect 113514 -1862 113546 -1626
rect 113782 -1862 113866 -1626
rect 114102 -1862 114134 -1626
rect 113514 -7654 114134 -1862
rect 117234 10894 117854 12559
rect 117234 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 117854 10894
rect 117234 10574 117854 10658
rect 117234 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 117854 10574
rect 117234 -2266 117854 10338
rect 117234 -2502 117266 -2266
rect 117502 -2502 117586 -2266
rect 117822 -2502 117854 -2266
rect 117234 -2586 117854 -2502
rect 117234 -2822 117266 -2586
rect 117502 -2822 117586 -2586
rect 117822 -2822 117854 -2586
rect 117234 -7654 117854 -2822
rect 145794 3454 146414 12559
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -7654 146414 -902
rect 149514 7174 150134 12559
rect 149514 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 150134 7174
rect 149514 6854 150134 6938
rect 149514 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 150134 6854
rect 149514 -1306 150134 6618
rect 149514 -1542 149546 -1306
rect 149782 -1542 149866 -1306
rect 150102 -1542 150134 -1306
rect 149514 -1626 150134 -1542
rect 149514 -1862 149546 -1626
rect 149782 -1862 149866 -1626
rect 150102 -1862 150134 -1626
rect 149514 -7654 150134 -1862
rect 153234 10894 153854 12559
rect 153234 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 153854 10894
rect 153234 10574 153854 10658
rect 153234 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 153854 10574
rect 153234 -2266 153854 10338
rect 153234 -2502 153266 -2266
rect 153502 -2502 153586 -2266
rect 153822 -2502 153854 -2266
rect 153234 -2586 153854 -2502
rect 153234 -2822 153266 -2586
rect 153502 -2822 153586 -2586
rect 153822 -2822 153854 -2586
rect 153234 -7654 153854 -2822
rect 181794 3454 182414 12559
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -7654 182414 -902
rect 185514 7174 186134 12068
rect 185514 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 186134 7174
rect 185514 6854 186134 6938
rect 185514 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 186134 6854
rect 185514 -1306 186134 6618
rect 185514 -1542 185546 -1306
rect 185782 -1542 185866 -1306
rect 186102 -1542 186134 -1306
rect 185514 -1626 186134 -1542
rect 185514 -1862 185546 -1626
rect 185782 -1862 185866 -1626
rect 186102 -1862 186134 -1626
rect 185514 -7654 186134 -1862
rect 189234 10894 189854 12559
rect 189234 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 189854 10894
rect 189234 10574 189854 10658
rect 189234 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 189854 10574
rect 189234 -2266 189854 10338
rect 189234 -2502 189266 -2266
rect 189502 -2502 189586 -2266
rect 189822 -2502 189854 -2266
rect 189234 -2586 189854 -2502
rect 189234 -2822 189266 -2586
rect 189502 -2822 189586 -2586
rect 189822 -2822 189854 -2586
rect 189234 -7654 189854 -2822
rect 217794 3454 218414 12559
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -7654 218414 -902
rect 221514 7174 222134 12559
rect 221514 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 222134 7174
rect 221514 6854 222134 6938
rect 221514 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 222134 6854
rect 221514 -1306 222134 6618
rect 221514 -1542 221546 -1306
rect 221782 -1542 221866 -1306
rect 222102 -1542 222134 -1306
rect 221514 -1626 222134 -1542
rect 221514 -1862 221546 -1626
rect 221782 -1862 221866 -1626
rect 222102 -1862 222134 -1626
rect 221514 -7654 222134 -1862
rect 225234 10894 225854 12559
rect 225234 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 225854 10894
rect 225234 10574 225854 10658
rect 225234 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 225854 10574
rect 225234 -2266 225854 10338
rect 225234 -2502 225266 -2266
rect 225502 -2502 225586 -2266
rect 225822 -2502 225854 -2266
rect 225234 -2586 225854 -2502
rect 225234 -2822 225266 -2586
rect 225502 -2822 225586 -2586
rect 225822 -2822 225854 -2586
rect 225234 -7654 225854 -2822
rect 253794 3454 254414 12559
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -7654 254414 -902
rect 257514 7174 258134 12559
rect 257514 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 258134 7174
rect 257514 6854 258134 6938
rect 257514 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 258134 6854
rect 257514 -1306 258134 6618
rect 257514 -1542 257546 -1306
rect 257782 -1542 257866 -1306
rect 258102 -1542 258134 -1306
rect 257514 -1626 258134 -1542
rect 257514 -1862 257546 -1626
rect 257782 -1862 257866 -1626
rect 258102 -1862 258134 -1626
rect 257514 -7654 258134 -1862
rect 261234 10894 261854 12559
rect 261234 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 261854 10894
rect 261234 10574 261854 10658
rect 261234 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 261854 10574
rect 261234 -2266 261854 10338
rect 261234 -2502 261266 -2266
rect 261502 -2502 261586 -2266
rect 261822 -2502 261854 -2266
rect 261234 -2586 261854 -2502
rect 261234 -2822 261266 -2586
rect 261502 -2822 261586 -2586
rect 261822 -2822 261854 -2586
rect 261234 -7654 261854 -2822
rect 289794 3454 290414 12559
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -7654 290414 -902
rect 293514 7174 294134 12559
rect 293514 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 294134 7174
rect 293514 6854 294134 6938
rect 293514 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 294134 6854
rect 293514 -1306 294134 6618
rect 293514 -1542 293546 -1306
rect 293782 -1542 293866 -1306
rect 294102 -1542 294134 -1306
rect 293514 -1626 294134 -1542
rect 293514 -1862 293546 -1626
rect 293782 -1862 293866 -1626
rect 294102 -1862 294134 -1626
rect 293514 -7654 294134 -1862
rect 297234 10894 297854 12559
rect 297234 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 297854 10894
rect 297234 10574 297854 10658
rect 297234 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 297854 10574
rect 297234 -2266 297854 10338
rect 297234 -2502 297266 -2266
rect 297502 -2502 297586 -2266
rect 297822 -2502 297854 -2266
rect 297234 -2586 297854 -2502
rect 297234 -2822 297266 -2586
rect 297502 -2822 297586 -2586
rect 297822 -2822 297854 -2586
rect 297234 -7654 297854 -2822
rect 325794 3454 326414 12559
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -7654 326414 -902
rect 329514 7174 330134 12559
rect 329514 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 330134 7174
rect 329514 6854 330134 6938
rect 329514 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 330134 6854
rect 329514 -1306 330134 6618
rect 329514 -1542 329546 -1306
rect 329782 -1542 329866 -1306
rect 330102 -1542 330134 -1306
rect 329514 -1626 330134 -1542
rect 329514 -1862 329546 -1626
rect 329782 -1862 329866 -1626
rect 330102 -1862 330134 -1626
rect 329514 -7654 330134 -1862
rect 333234 10894 333854 12559
rect 333234 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 333854 10894
rect 333234 10574 333854 10658
rect 333234 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 333854 10574
rect 333234 -2266 333854 10338
rect 333234 -2502 333266 -2266
rect 333502 -2502 333586 -2266
rect 333822 -2502 333854 -2266
rect 333234 -2586 333854 -2502
rect 333234 -2822 333266 -2586
rect 333502 -2822 333586 -2586
rect 333822 -2822 333854 -2586
rect 333234 -7654 333854 -2822
rect 361794 3454 362414 12559
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -7654 362414 -902
rect 365514 7174 366134 12559
rect 365514 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 366134 7174
rect 365514 6854 366134 6938
rect 365514 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 366134 6854
rect 365514 -1306 366134 6618
rect 365514 -1542 365546 -1306
rect 365782 -1542 365866 -1306
rect 366102 -1542 366134 -1306
rect 365514 -1626 366134 -1542
rect 365514 -1862 365546 -1626
rect 365782 -1862 365866 -1626
rect 366102 -1862 366134 -1626
rect 365514 -7654 366134 -1862
rect 369234 10894 369854 12068
rect 369234 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 369854 10894
rect 369234 10574 369854 10658
rect 369234 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 369854 10574
rect 369234 -2266 369854 10338
rect 369234 -2502 369266 -2266
rect 369502 -2502 369586 -2266
rect 369822 -2502 369854 -2266
rect 369234 -2586 369854 -2502
rect 369234 -2822 369266 -2586
rect 369502 -2822 369586 -2586
rect 369822 -2822 369854 -2586
rect 369234 -7654 369854 -2822
rect 397794 3454 398414 12559
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -7654 398414 -902
rect 401514 7174 402134 12559
rect 401514 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 402134 7174
rect 401514 6854 402134 6938
rect 401514 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 402134 6854
rect 401514 -1306 402134 6618
rect 401514 -1542 401546 -1306
rect 401782 -1542 401866 -1306
rect 402102 -1542 402134 -1306
rect 401514 -1626 402134 -1542
rect 401514 -1862 401546 -1626
rect 401782 -1862 401866 -1626
rect 402102 -1862 402134 -1626
rect 401514 -7654 402134 -1862
rect 405234 10894 405854 12559
rect 405234 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 405854 10894
rect 405234 10574 405854 10658
rect 405234 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 405854 10574
rect 405234 -2266 405854 10338
rect 405234 -2502 405266 -2266
rect 405502 -2502 405586 -2266
rect 405822 -2502 405854 -2266
rect 405234 -2586 405854 -2502
rect 405234 -2822 405266 -2586
rect 405502 -2822 405586 -2586
rect 405822 -2822 405854 -2586
rect 405234 -7654 405854 -2822
rect 433794 3454 434414 12559
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -7654 434414 -902
rect 437514 7174 438134 12559
rect 437514 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 438134 7174
rect 437514 6854 438134 6938
rect 437514 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 438134 6854
rect 437514 -1306 438134 6618
rect 437514 -1542 437546 -1306
rect 437782 -1542 437866 -1306
rect 438102 -1542 438134 -1306
rect 437514 -1626 438134 -1542
rect 437514 -1862 437546 -1626
rect 437782 -1862 437866 -1626
rect 438102 -1862 438134 -1626
rect 437514 -7654 438134 -1862
rect 441234 10894 441854 12559
rect 441234 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 441854 10894
rect 441234 10574 441854 10658
rect 441234 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 441854 10574
rect 441234 -2266 441854 10338
rect 441234 -2502 441266 -2266
rect 441502 -2502 441586 -2266
rect 441822 -2502 441854 -2266
rect 441234 -2586 441854 -2502
rect 441234 -2822 441266 -2586
rect 441502 -2822 441586 -2586
rect 441822 -2822 441854 -2586
rect 441234 -7654 441854 -2822
rect 469794 3454 470414 12559
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -7654 470414 -902
rect 473514 7174 474134 12559
rect 473514 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 474134 7174
rect 473514 6854 474134 6938
rect 473514 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 474134 6854
rect 473514 -1306 474134 6618
rect 473514 -1542 473546 -1306
rect 473782 -1542 473866 -1306
rect 474102 -1542 474134 -1306
rect 473514 -1626 474134 -1542
rect 473514 -1862 473546 -1626
rect 473782 -1862 473866 -1626
rect 474102 -1862 474134 -1626
rect 473514 -7654 474134 -1862
rect 477234 10894 477854 12068
rect 477234 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 477854 10894
rect 477234 10574 477854 10658
rect 477234 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 477854 10574
rect 477234 -2266 477854 10338
rect 477234 -2502 477266 -2266
rect 477502 -2502 477586 -2266
rect 477822 -2502 477854 -2266
rect 477234 -2586 477854 -2502
rect 477234 -2822 477266 -2586
rect 477502 -2822 477586 -2586
rect 477822 -2822 477854 -2586
rect 477234 -7654 477854 -2822
rect 505794 3454 506414 12559
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -7654 506414 -902
rect 509514 7174 510134 12559
rect 509514 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 510134 7174
rect 509514 6854 510134 6938
rect 509514 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 510134 6854
rect 509514 -1306 510134 6618
rect 509514 -1542 509546 -1306
rect 509782 -1542 509866 -1306
rect 510102 -1542 510134 -1306
rect 509514 -1626 510134 -1542
rect 509514 -1862 509546 -1626
rect 509782 -1862 509866 -1626
rect 510102 -1862 510134 -1626
rect 509514 -7654 510134 -1862
rect 513234 10894 513854 12559
rect 513234 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 513854 10894
rect 513234 10574 513854 10658
rect 513234 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 513854 10574
rect 513234 -2266 513854 10338
rect 513234 -2502 513266 -2266
rect 513502 -2502 513586 -2266
rect 513822 -2502 513854 -2266
rect 513234 -2586 513854 -2502
rect 513234 -2822 513266 -2586
rect 513502 -2822 513586 -2586
rect 513822 -2822 513854 -2586
rect 513234 -7654 513854 -2822
rect 541794 3454 542414 12559
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -7654 542414 -902
rect 545514 7174 546134 12559
rect 545514 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 546134 7174
rect 545514 6854 546134 6938
rect 545514 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 546134 6854
rect 545514 -1306 546134 6618
rect 545514 -1542 545546 -1306
rect 545782 -1542 545866 -1306
rect 546102 -1542 546134 -1306
rect 545514 -1626 546134 -1542
rect 545514 -1862 545546 -1626
rect 545782 -1862 545866 -1626
rect 546102 -1862 546134 -1626
rect 545514 -7654 546134 -1862
rect 549234 10894 549854 12559
rect 549234 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 549854 10894
rect 549234 10574 549854 10658
rect 549234 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 549854 10574
rect 549234 -2266 549854 10338
rect 549234 -2502 549266 -2266
rect 549502 -2502 549586 -2266
rect 549822 -2502 549854 -2266
rect 549234 -2586 549854 -2502
rect 549234 -2822 549266 -2586
rect 549502 -2822 549586 -2586
rect 549822 -2822 549854 -2586
rect 549234 -7654 549854 -2822
rect 567834 -7066 568454 28938
rect 567834 -7302 567866 -7066
rect 568102 -7302 568186 -7066
rect 568422 -7302 568454 -7066
rect 567834 -7386 568454 -7302
rect 567834 -7622 567866 -7386
rect 568102 -7622 568186 -7386
rect 568422 -7622 568454 -7386
rect 567834 -7654 568454 -7622
rect 577794 704838 578414 711590
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -7654 578414 -902
rect 581514 705798 582134 711590
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 581514 705562 581546 705798
rect 581782 705562 581866 705798
rect 582102 705562 582134 705798
rect 581514 705478 582134 705562
rect 581514 705242 581546 705478
rect 581782 705242 581866 705478
rect 582102 705242 582134 705478
rect 581514 691174 582134 705242
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 581514 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 582134 691174
rect 581514 690854 582134 690938
rect 581514 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 582134 690854
rect 581514 655174 582134 690618
rect 581514 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 582134 655174
rect 581514 654854 582134 654938
rect 581514 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 582134 654854
rect 581514 619174 582134 654618
rect 581514 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 582134 619174
rect 581514 618854 582134 618938
rect 581514 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 582134 618854
rect 581514 583174 582134 618618
rect 581514 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 582134 583174
rect 581514 582854 582134 582938
rect 581514 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 582134 582854
rect 581514 547174 582134 582618
rect 581514 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 582134 547174
rect 581514 546854 582134 546938
rect 581514 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 582134 546854
rect 581514 511174 582134 546618
rect 581514 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 582134 511174
rect 581514 510854 582134 510938
rect 581514 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 582134 510854
rect 581514 475174 582134 510618
rect 581514 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 582134 475174
rect 581514 474854 582134 474938
rect 581514 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 582134 474854
rect 581514 439174 582134 474618
rect 581514 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 582134 439174
rect 581514 438854 582134 438938
rect 581514 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 582134 438854
rect 581514 403174 582134 438618
rect 581514 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 582134 403174
rect 581514 402854 582134 402938
rect 581514 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 582134 402854
rect 581514 367174 582134 402618
rect 581514 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 582134 367174
rect 581514 366854 582134 366938
rect 581514 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 582134 366854
rect 581514 331174 582134 366618
rect 581514 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 582134 331174
rect 581514 330854 582134 330938
rect 581514 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 582134 330854
rect 581514 295174 582134 330618
rect 581514 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 582134 295174
rect 581514 294854 582134 294938
rect 581514 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 582134 294854
rect 581514 259174 582134 294618
rect 581514 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 582134 259174
rect 581514 258854 582134 258938
rect 581514 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 582134 258854
rect 581514 223174 582134 258618
rect 581514 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 582134 223174
rect 581514 222854 582134 222938
rect 581514 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 582134 222854
rect 581514 187174 582134 222618
rect 581514 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 582134 187174
rect 581514 186854 582134 186938
rect 581514 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 582134 186854
rect 581514 151174 582134 186618
rect 581514 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 582134 151174
rect 581514 150854 582134 150938
rect 581514 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 582134 150854
rect 581514 115174 582134 150618
rect 581514 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 582134 115174
rect 581514 114854 582134 114938
rect 581514 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 582134 114854
rect 581514 79174 582134 114618
rect 581514 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 582134 79174
rect 581514 78854 582134 78938
rect 581514 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 582134 78854
rect 581514 43174 582134 78618
rect 581514 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 582134 43174
rect 581514 42854 582134 42938
rect 581514 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 582134 42854
rect 581514 7174 582134 42618
rect 581514 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 582134 7174
rect 581514 6854 582134 6938
rect 581514 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 582134 6854
rect 581514 -1306 582134 6618
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 691174 586890 705242
rect 586270 690938 586302 691174
rect 586538 690938 586622 691174
rect 586858 690938 586890 691174
rect 586270 690854 586890 690938
rect 586270 690618 586302 690854
rect 586538 690618 586622 690854
rect 586858 690618 586890 690854
rect 586270 655174 586890 690618
rect 586270 654938 586302 655174
rect 586538 654938 586622 655174
rect 586858 654938 586890 655174
rect 586270 654854 586890 654938
rect 586270 654618 586302 654854
rect 586538 654618 586622 654854
rect 586858 654618 586890 654854
rect 586270 619174 586890 654618
rect 586270 618938 586302 619174
rect 586538 618938 586622 619174
rect 586858 618938 586890 619174
rect 586270 618854 586890 618938
rect 586270 618618 586302 618854
rect 586538 618618 586622 618854
rect 586858 618618 586890 618854
rect 586270 583174 586890 618618
rect 586270 582938 586302 583174
rect 586538 582938 586622 583174
rect 586858 582938 586890 583174
rect 586270 582854 586890 582938
rect 586270 582618 586302 582854
rect 586538 582618 586622 582854
rect 586858 582618 586890 582854
rect 586270 547174 586890 582618
rect 586270 546938 586302 547174
rect 586538 546938 586622 547174
rect 586858 546938 586890 547174
rect 586270 546854 586890 546938
rect 586270 546618 586302 546854
rect 586538 546618 586622 546854
rect 586858 546618 586890 546854
rect 586270 511174 586890 546618
rect 586270 510938 586302 511174
rect 586538 510938 586622 511174
rect 586858 510938 586890 511174
rect 586270 510854 586890 510938
rect 586270 510618 586302 510854
rect 586538 510618 586622 510854
rect 586858 510618 586890 510854
rect 586270 475174 586890 510618
rect 586270 474938 586302 475174
rect 586538 474938 586622 475174
rect 586858 474938 586890 475174
rect 586270 474854 586890 474938
rect 586270 474618 586302 474854
rect 586538 474618 586622 474854
rect 586858 474618 586890 474854
rect 586270 439174 586890 474618
rect 586270 438938 586302 439174
rect 586538 438938 586622 439174
rect 586858 438938 586890 439174
rect 586270 438854 586890 438938
rect 586270 438618 586302 438854
rect 586538 438618 586622 438854
rect 586858 438618 586890 438854
rect 586270 403174 586890 438618
rect 586270 402938 586302 403174
rect 586538 402938 586622 403174
rect 586858 402938 586890 403174
rect 586270 402854 586890 402938
rect 586270 402618 586302 402854
rect 586538 402618 586622 402854
rect 586858 402618 586890 402854
rect 586270 367174 586890 402618
rect 586270 366938 586302 367174
rect 586538 366938 586622 367174
rect 586858 366938 586890 367174
rect 586270 366854 586890 366938
rect 586270 366618 586302 366854
rect 586538 366618 586622 366854
rect 586858 366618 586890 366854
rect 586270 331174 586890 366618
rect 586270 330938 586302 331174
rect 586538 330938 586622 331174
rect 586858 330938 586890 331174
rect 586270 330854 586890 330938
rect 586270 330618 586302 330854
rect 586538 330618 586622 330854
rect 586858 330618 586890 330854
rect 586270 295174 586890 330618
rect 586270 294938 586302 295174
rect 586538 294938 586622 295174
rect 586858 294938 586890 295174
rect 586270 294854 586890 294938
rect 586270 294618 586302 294854
rect 586538 294618 586622 294854
rect 586858 294618 586890 294854
rect 586270 259174 586890 294618
rect 586270 258938 586302 259174
rect 586538 258938 586622 259174
rect 586858 258938 586890 259174
rect 586270 258854 586890 258938
rect 586270 258618 586302 258854
rect 586538 258618 586622 258854
rect 586858 258618 586890 258854
rect 586270 223174 586890 258618
rect 586270 222938 586302 223174
rect 586538 222938 586622 223174
rect 586858 222938 586890 223174
rect 586270 222854 586890 222938
rect 586270 222618 586302 222854
rect 586538 222618 586622 222854
rect 586858 222618 586890 222854
rect 586270 187174 586890 222618
rect 586270 186938 586302 187174
rect 586538 186938 586622 187174
rect 586858 186938 586890 187174
rect 586270 186854 586890 186938
rect 586270 186618 586302 186854
rect 586538 186618 586622 186854
rect 586858 186618 586890 186854
rect 586270 151174 586890 186618
rect 586270 150938 586302 151174
rect 586538 150938 586622 151174
rect 586858 150938 586890 151174
rect 586270 150854 586890 150938
rect 586270 150618 586302 150854
rect 586538 150618 586622 150854
rect 586858 150618 586890 150854
rect 586270 115174 586890 150618
rect 586270 114938 586302 115174
rect 586538 114938 586622 115174
rect 586858 114938 586890 115174
rect 586270 114854 586890 114938
rect 586270 114618 586302 114854
rect 586538 114618 586622 114854
rect 586858 114618 586890 114854
rect 586270 79174 586890 114618
rect 586270 78938 586302 79174
rect 586538 78938 586622 79174
rect 586858 78938 586890 79174
rect 586270 78854 586890 78938
rect 586270 78618 586302 78854
rect 586538 78618 586622 78854
rect 586858 78618 586890 78854
rect 586270 43174 586890 78618
rect 586270 42938 586302 43174
rect 586538 42938 586622 43174
rect 586858 42938 586890 43174
rect 586270 42854 586890 42938
rect 586270 42618 586302 42854
rect 586538 42618 586622 42854
rect 586858 42618 586890 42854
rect 586270 7174 586890 42618
rect 586270 6938 586302 7174
rect 586538 6938 586622 7174
rect 586858 6938 586890 7174
rect 586270 6854 586890 6938
rect 586270 6618 586302 6854
rect 586538 6618 586622 6854
rect 586858 6618 586890 6854
rect 581514 -1542 581546 -1306
rect 581782 -1542 581866 -1306
rect 582102 -1542 582134 -1306
rect 581514 -1626 582134 -1542
rect 581514 -1862 581546 -1626
rect 581782 -1862 581866 -1626
rect 582102 -1862 582134 -1626
rect 581514 -7654 582134 -1862
rect 586270 -1306 586890 6618
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 694894 587850 706202
rect 587230 694658 587262 694894
rect 587498 694658 587582 694894
rect 587818 694658 587850 694894
rect 587230 694574 587850 694658
rect 587230 694338 587262 694574
rect 587498 694338 587582 694574
rect 587818 694338 587850 694574
rect 587230 658894 587850 694338
rect 587230 658658 587262 658894
rect 587498 658658 587582 658894
rect 587818 658658 587850 658894
rect 587230 658574 587850 658658
rect 587230 658338 587262 658574
rect 587498 658338 587582 658574
rect 587818 658338 587850 658574
rect 587230 622894 587850 658338
rect 587230 622658 587262 622894
rect 587498 622658 587582 622894
rect 587818 622658 587850 622894
rect 587230 622574 587850 622658
rect 587230 622338 587262 622574
rect 587498 622338 587582 622574
rect 587818 622338 587850 622574
rect 587230 586894 587850 622338
rect 587230 586658 587262 586894
rect 587498 586658 587582 586894
rect 587818 586658 587850 586894
rect 587230 586574 587850 586658
rect 587230 586338 587262 586574
rect 587498 586338 587582 586574
rect 587818 586338 587850 586574
rect 587230 550894 587850 586338
rect 587230 550658 587262 550894
rect 587498 550658 587582 550894
rect 587818 550658 587850 550894
rect 587230 550574 587850 550658
rect 587230 550338 587262 550574
rect 587498 550338 587582 550574
rect 587818 550338 587850 550574
rect 587230 514894 587850 550338
rect 587230 514658 587262 514894
rect 587498 514658 587582 514894
rect 587818 514658 587850 514894
rect 587230 514574 587850 514658
rect 587230 514338 587262 514574
rect 587498 514338 587582 514574
rect 587818 514338 587850 514574
rect 587230 478894 587850 514338
rect 587230 478658 587262 478894
rect 587498 478658 587582 478894
rect 587818 478658 587850 478894
rect 587230 478574 587850 478658
rect 587230 478338 587262 478574
rect 587498 478338 587582 478574
rect 587818 478338 587850 478574
rect 587230 442894 587850 478338
rect 587230 442658 587262 442894
rect 587498 442658 587582 442894
rect 587818 442658 587850 442894
rect 587230 442574 587850 442658
rect 587230 442338 587262 442574
rect 587498 442338 587582 442574
rect 587818 442338 587850 442574
rect 587230 406894 587850 442338
rect 587230 406658 587262 406894
rect 587498 406658 587582 406894
rect 587818 406658 587850 406894
rect 587230 406574 587850 406658
rect 587230 406338 587262 406574
rect 587498 406338 587582 406574
rect 587818 406338 587850 406574
rect 587230 370894 587850 406338
rect 587230 370658 587262 370894
rect 587498 370658 587582 370894
rect 587818 370658 587850 370894
rect 587230 370574 587850 370658
rect 587230 370338 587262 370574
rect 587498 370338 587582 370574
rect 587818 370338 587850 370574
rect 587230 334894 587850 370338
rect 587230 334658 587262 334894
rect 587498 334658 587582 334894
rect 587818 334658 587850 334894
rect 587230 334574 587850 334658
rect 587230 334338 587262 334574
rect 587498 334338 587582 334574
rect 587818 334338 587850 334574
rect 587230 298894 587850 334338
rect 587230 298658 587262 298894
rect 587498 298658 587582 298894
rect 587818 298658 587850 298894
rect 587230 298574 587850 298658
rect 587230 298338 587262 298574
rect 587498 298338 587582 298574
rect 587818 298338 587850 298574
rect 587230 262894 587850 298338
rect 587230 262658 587262 262894
rect 587498 262658 587582 262894
rect 587818 262658 587850 262894
rect 587230 262574 587850 262658
rect 587230 262338 587262 262574
rect 587498 262338 587582 262574
rect 587818 262338 587850 262574
rect 587230 226894 587850 262338
rect 587230 226658 587262 226894
rect 587498 226658 587582 226894
rect 587818 226658 587850 226894
rect 587230 226574 587850 226658
rect 587230 226338 587262 226574
rect 587498 226338 587582 226574
rect 587818 226338 587850 226574
rect 587230 190894 587850 226338
rect 587230 190658 587262 190894
rect 587498 190658 587582 190894
rect 587818 190658 587850 190894
rect 587230 190574 587850 190658
rect 587230 190338 587262 190574
rect 587498 190338 587582 190574
rect 587818 190338 587850 190574
rect 587230 154894 587850 190338
rect 587230 154658 587262 154894
rect 587498 154658 587582 154894
rect 587818 154658 587850 154894
rect 587230 154574 587850 154658
rect 587230 154338 587262 154574
rect 587498 154338 587582 154574
rect 587818 154338 587850 154574
rect 587230 118894 587850 154338
rect 587230 118658 587262 118894
rect 587498 118658 587582 118894
rect 587818 118658 587850 118894
rect 587230 118574 587850 118658
rect 587230 118338 587262 118574
rect 587498 118338 587582 118574
rect 587818 118338 587850 118574
rect 587230 82894 587850 118338
rect 587230 82658 587262 82894
rect 587498 82658 587582 82894
rect 587818 82658 587850 82894
rect 587230 82574 587850 82658
rect 587230 82338 587262 82574
rect 587498 82338 587582 82574
rect 587818 82338 587850 82574
rect 587230 46894 587850 82338
rect 587230 46658 587262 46894
rect 587498 46658 587582 46894
rect 587818 46658 587850 46894
rect 587230 46574 587850 46658
rect 587230 46338 587262 46574
rect 587498 46338 587582 46574
rect 587818 46338 587850 46574
rect 587230 10894 587850 46338
rect 587230 10658 587262 10894
rect 587498 10658 587582 10894
rect 587818 10658 587850 10894
rect 587230 10574 587850 10658
rect 587230 10338 587262 10574
rect 587498 10338 587582 10574
rect 587818 10338 587850 10574
rect 587230 -2266 587850 10338
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 698614 588810 707162
rect 588190 698378 588222 698614
rect 588458 698378 588542 698614
rect 588778 698378 588810 698614
rect 588190 698294 588810 698378
rect 588190 698058 588222 698294
rect 588458 698058 588542 698294
rect 588778 698058 588810 698294
rect 588190 662614 588810 698058
rect 588190 662378 588222 662614
rect 588458 662378 588542 662614
rect 588778 662378 588810 662614
rect 588190 662294 588810 662378
rect 588190 662058 588222 662294
rect 588458 662058 588542 662294
rect 588778 662058 588810 662294
rect 588190 626614 588810 662058
rect 588190 626378 588222 626614
rect 588458 626378 588542 626614
rect 588778 626378 588810 626614
rect 588190 626294 588810 626378
rect 588190 626058 588222 626294
rect 588458 626058 588542 626294
rect 588778 626058 588810 626294
rect 588190 590614 588810 626058
rect 588190 590378 588222 590614
rect 588458 590378 588542 590614
rect 588778 590378 588810 590614
rect 588190 590294 588810 590378
rect 588190 590058 588222 590294
rect 588458 590058 588542 590294
rect 588778 590058 588810 590294
rect 588190 554614 588810 590058
rect 588190 554378 588222 554614
rect 588458 554378 588542 554614
rect 588778 554378 588810 554614
rect 588190 554294 588810 554378
rect 588190 554058 588222 554294
rect 588458 554058 588542 554294
rect 588778 554058 588810 554294
rect 588190 518614 588810 554058
rect 588190 518378 588222 518614
rect 588458 518378 588542 518614
rect 588778 518378 588810 518614
rect 588190 518294 588810 518378
rect 588190 518058 588222 518294
rect 588458 518058 588542 518294
rect 588778 518058 588810 518294
rect 588190 482614 588810 518058
rect 588190 482378 588222 482614
rect 588458 482378 588542 482614
rect 588778 482378 588810 482614
rect 588190 482294 588810 482378
rect 588190 482058 588222 482294
rect 588458 482058 588542 482294
rect 588778 482058 588810 482294
rect 588190 446614 588810 482058
rect 588190 446378 588222 446614
rect 588458 446378 588542 446614
rect 588778 446378 588810 446614
rect 588190 446294 588810 446378
rect 588190 446058 588222 446294
rect 588458 446058 588542 446294
rect 588778 446058 588810 446294
rect 588190 410614 588810 446058
rect 588190 410378 588222 410614
rect 588458 410378 588542 410614
rect 588778 410378 588810 410614
rect 588190 410294 588810 410378
rect 588190 410058 588222 410294
rect 588458 410058 588542 410294
rect 588778 410058 588810 410294
rect 588190 374614 588810 410058
rect 588190 374378 588222 374614
rect 588458 374378 588542 374614
rect 588778 374378 588810 374614
rect 588190 374294 588810 374378
rect 588190 374058 588222 374294
rect 588458 374058 588542 374294
rect 588778 374058 588810 374294
rect 588190 338614 588810 374058
rect 588190 338378 588222 338614
rect 588458 338378 588542 338614
rect 588778 338378 588810 338614
rect 588190 338294 588810 338378
rect 588190 338058 588222 338294
rect 588458 338058 588542 338294
rect 588778 338058 588810 338294
rect 588190 302614 588810 338058
rect 588190 302378 588222 302614
rect 588458 302378 588542 302614
rect 588778 302378 588810 302614
rect 588190 302294 588810 302378
rect 588190 302058 588222 302294
rect 588458 302058 588542 302294
rect 588778 302058 588810 302294
rect 588190 266614 588810 302058
rect 588190 266378 588222 266614
rect 588458 266378 588542 266614
rect 588778 266378 588810 266614
rect 588190 266294 588810 266378
rect 588190 266058 588222 266294
rect 588458 266058 588542 266294
rect 588778 266058 588810 266294
rect 588190 230614 588810 266058
rect 588190 230378 588222 230614
rect 588458 230378 588542 230614
rect 588778 230378 588810 230614
rect 588190 230294 588810 230378
rect 588190 230058 588222 230294
rect 588458 230058 588542 230294
rect 588778 230058 588810 230294
rect 588190 194614 588810 230058
rect 588190 194378 588222 194614
rect 588458 194378 588542 194614
rect 588778 194378 588810 194614
rect 588190 194294 588810 194378
rect 588190 194058 588222 194294
rect 588458 194058 588542 194294
rect 588778 194058 588810 194294
rect 588190 158614 588810 194058
rect 588190 158378 588222 158614
rect 588458 158378 588542 158614
rect 588778 158378 588810 158614
rect 588190 158294 588810 158378
rect 588190 158058 588222 158294
rect 588458 158058 588542 158294
rect 588778 158058 588810 158294
rect 588190 122614 588810 158058
rect 588190 122378 588222 122614
rect 588458 122378 588542 122614
rect 588778 122378 588810 122614
rect 588190 122294 588810 122378
rect 588190 122058 588222 122294
rect 588458 122058 588542 122294
rect 588778 122058 588810 122294
rect 588190 86614 588810 122058
rect 588190 86378 588222 86614
rect 588458 86378 588542 86614
rect 588778 86378 588810 86614
rect 588190 86294 588810 86378
rect 588190 86058 588222 86294
rect 588458 86058 588542 86294
rect 588778 86058 588810 86294
rect 588190 50614 588810 86058
rect 588190 50378 588222 50614
rect 588458 50378 588542 50614
rect 588778 50378 588810 50614
rect 588190 50294 588810 50378
rect 588190 50058 588222 50294
rect 588458 50058 588542 50294
rect 588778 50058 588810 50294
rect 588190 14614 588810 50058
rect 588190 14378 588222 14614
rect 588458 14378 588542 14614
rect 588778 14378 588810 14614
rect 588190 14294 588810 14378
rect 588190 14058 588222 14294
rect 588458 14058 588542 14294
rect 588778 14058 588810 14294
rect 588190 -3226 588810 14058
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 666334 589770 708122
rect 589150 666098 589182 666334
rect 589418 666098 589502 666334
rect 589738 666098 589770 666334
rect 589150 666014 589770 666098
rect 589150 665778 589182 666014
rect 589418 665778 589502 666014
rect 589738 665778 589770 666014
rect 589150 630334 589770 665778
rect 589150 630098 589182 630334
rect 589418 630098 589502 630334
rect 589738 630098 589770 630334
rect 589150 630014 589770 630098
rect 589150 629778 589182 630014
rect 589418 629778 589502 630014
rect 589738 629778 589770 630014
rect 589150 594334 589770 629778
rect 589150 594098 589182 594334
rect 589418 594098 589502 594334
rect 589738 594098 589770 594334
rect 589150 594014 589770 594098
rect 589150 593778 589182 594014
rect 589418 593778 589502 594014
rect 589738 593778 589770 594014
rect 589150 558334 589770 593778
rect 589150 558098 589182 558334
rect 589418 558098 589502 558334
rect 589738 558098 589770 558334
rect 589150 558014 589770 558098
rect 589150 557778 589182 558014
rect 589418 557778 589502 558014
rect 589738 557778 589770 558014
rect 589150 522334 589770 557778
rect 589150 522098 589182 522334
rect 589418 522098 589502 522334
rect 589738 522098 589770 522334
rect 589150 522014 589770 522098
rect 589150 521778 589182 522014
rect 589418 521778 589502 522014
rect 589738 521778 589770 522014
rect 589150 486334 589770 521778
rect 589150 486098 589182 486334
rect 589418 486098 589502 486334
rect 589738 486098 589770 486334
rect 589150 486014 589770 486098
rect 589150 485778 589182 486014
rect 589418 485778 589502 486014
rect 589738 485778 589770 486014
rect 589150 450334 589770 485778
rect 589150 450098 589182 450334
rect 589418 450098 589502 450334
rect 589738 450098 589770 450334
rect 589150 450014 589770 450098
rect 589150 449778 589182 450014
rect 589418 449778 589502 450014
rect 589738 449778 589770 450014
rect 589150 414334 589770 449778
rect 589150 414098 589182 414334
rect 589418 414098 589502 414334
rect 589738 414098 589770 414334
rect 589150 414014 589770 414098
rect 589150 413778 589182 414014
rect 589418 413778 589502 414014
rect 589738 413778 589770 414014
rect 589150 378334 589770 413778
rect 589150 378098 589182 378334
rect 589418 378098 589502 378334
rect 589738 378098 589770 378334
rect 589150 378014 589770 378098
rect 589150 377778 589182 378014
rect 589418 377778 589502 378014
rect 589738 377778 589770 378014
rect 589150 342334 589770 377778
rect 589150 342098 589182 342334
rect 589418 342098 589502 342334
rect 589738 342098 589770 342334
rect 589150 342014 589770 342098
rect 589150 341778 589182 342014
rect 589418 341778 589502 342014
rect 589738 341778 589770 342014
rect 589150 306334 589770 341778
rect 589150 306098 589182 306334
rect 589418 306098 589502 306334
rect 589738 306098 589770 306334
rect 589150 306014 589770 306098
rect 589150 305778 589182 306014
rect 589418 305778 589502 306014
rect 589738 305778 589770 306014
rect 589150 270334 589770 305778
rect 589150 270098 589182 270334
rect 589418 270098 589502 270334
rect 589738 270098 589770 270334
rect 589150 270014 589770 270098
rect 589150 269778 589182 270014
rect 589418 269778 589502 270014
rect 589738 269778 589770 270014
rect 589150 234334 589770 269778
rect 589150 234098 589182 234334
rect 589418 234098 589502 234334
rect 589738 234098 589770 234334
rect 589150 234014 589770 234098
rect 589150 233778 589182 234014
rect 589418 233778 589502 234014
rect 589738 233778 589770 234014
rect 589150 198334 589770 233778
rect 589150 198098 589182 198334
rect 589418 198098 589502 198334
rect 589738 198098 589770 198334
rect 589150 198014 589770 198098
rect 589150 197778 589182 198014
rect 589418 197778 589502 198014
rect 589738 197778 589770 198014
rect 589150 162334 589770 197778
rect 589150 162098 589182 162334
rect 589418 162098 589502 162334
rect 589738 162098 589770 162334
rect 589150 162014 589770 162098
rect 589150 161778 589182 162014
rect 589418 161778 589502 162014
rect 589738 161778 589770 162014
rect 589150 126334 589770 161778
rect 589150 126098 589182 126334
rect 589418 126098 589502 126334
rect 589738 126098 589770 126334
rect 589150 126014 589770 126098
rect 589150 125778 589182 126014
rect 589418 125778 589502 126014
rect 589738 125778 589770 126014
rect 589150 90334 589770 125778
rect 589150 90098 589182 90334
rect 589418 90098 589502 90334
rect 589738 90098 589770 90334
rect 589150 90014 589770 90098
rect 589150 89778 589182 90014
rect 589418 89778 589502 90014
rect 589738 89778 589770 90014
rect 589150 54334 589770 89778
rect 589150 54098 589182 54334
rect 589418 54098 589502 54334
rect 589738 54098 589770 54334
rect 589150 54014 589770 54098
rect 589150 53778 589182 54014
rect 589418 53778 589502 54014
rect 589738 53778 589770 54014
rect 589150 18334 589770 53778
rect 589150 18098 589182 18334
rect 589418 18098 589502 18334
rect 589738 18098 589770 18334
rect 589150 18014 589770 18098
rect 589150 17778 589182 18014
rect 589418 17778 589502 18014
rect 589738 17778 589770 18014
rect 589150 -4186 589770 17778
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 670054 590730 709082
rect 590110 669818 590142 670054
rect 590378 669818 590462 670054
rect 590698 669818 590730 670054
rect 590110 669734 590730 669818
rect 590110 669498 590142 669734
rect 590378 669498 590462 669734
rect 590698 669498 590730 669734
rect 590110 634054 590730 669498
rect 590110 633818 590142 634054
rect 590378 633818 590462 634054
rect 590698 633818 590730 634054
rect 590110 633734 590730 633818
rect 590110 633498 590142 633734
rect 590378 633498 590462 633734
rect 590698 633498 590730 633734
rect 590110 598054 590730 633498
rect 590110 597818 590142 598054
rect 590378 597818 590462 598054
rect 590698 597818 590730 598054
rect 590110 597734 590730 597818
rect 590110 597498 590142 597734
rect 590378 597498 590462 597734
rect 590698 597498 590730 597734
rect 590110 562054 590730 597498
rect 590110 561818 590142 562054
rect 590378 561818 590462 562054
rect 590698 561818 590730 562054
rect 590110 561734 590730 561818
rect 590110 561498 590142 561734
rect 590378 561498 590462 561734
rect 590698 561498 590730 561734
rect 590110 526054 590730 561498
rect 590110 525818 590142 526054
rect 590378 525818 590462 526054
rect 590698 525818 590730 526054
rect 590110 525734 590730 525818
rect 590110 525498 590142 525734
rect 590378 525498 590462 525734
rect 590698 525498 590730 525734
rect 590110 490054 590730 525498
rect 590110 489818 590142 490054
rect 590378 489818 590462 490054
rect 590698 489818 590730 490054
rect 590110 489734 590730 489818
rect 590110 489498 590142 489734
rect 590378 489498 590462 489734
rect 590698 489498 590730 489734
rect 590110 454054 590730 489498
rect 590110 453818 590142 454054
rect 590378 453818 590462 454054
rect 590698 453818 590730 454054
rect 590110 453734 590730 453818
rect 590110 453498 590142 453734
rect 590378 453498 590462 453734
rect 590698 453498 590730 453734
rect 590110 418054 590730 453498
rect 590110 417818 590142 418054
rect 590378 417818 590462 418054
rect 590698 417818 590730 418054
rect 590110 417734 590730 417818
rect 590110 417498 590142 417734
rect 590378 417498 590462 417734
rect 590698 417498 590730 417734
rect 590110 382054 590730 417498
rect 590110 381818 590142 382054
rect 590378 381818 590462 382054
rect 590698 381818 590730 382054
rect 590110 381734 590730 381818
rect 590110 381498 590142 381734
rect 590378 381498 590462 381734
rect 590698 381498 590730 381734
rect 590110 346054 590730 381498
rect 590110 345818 590142 346054
rect 590378 345818 590462 346054
rect 590698 345818 590730 346054
rect 590110 345734 590730 345818
rect 590110 345498 590142 345734
rect 590378 345498 590462 345734
rect 590698 345498 590730 345734
rect 590110 310054 590730 345498
rect 590110 309818 590142 310054
rect 590378 309818 590462 310054
rect 590698 309818 590730 310054
rect 590110 309734 590730 309818
rect 590110 309498 590142 309734
rect 590378 309498 590462 309734
rect 590698 309498 590730 309734
rect 590110 274054 590730 309498
rect 590110 273818 590142 274054
rect 590378 273818 590462 274054
rect 590698 273818 590730 274054
rect 590110 273734 590730 273818
rect 590110 273498 590142 273734
rect 590378 273498 590462 273734
rect 590698 273498 590730 273734
rect 590110 238054 590730 273498
rect 590110 237818 590142 238054
rect 590378 237818 590462 238054
rect 590698 237818 590730 238054
rect 590110 237734 590730 237818
rect 590110 237498 590142 237734
rect 590378 237498 590462 237734
rect 590698 237498 590730 237734
rect 590110 202054 590730 237498
rect 590110 201818 590142 202054
rect 590378 201818 590462 202054
rect 590698 201818 590730 202054
rect 590110 201734 590730 201818
rect 590110 201498 590142 201734
rect 590378 201498 590462 201734
rect 590698 201498 590730 201734
rect 590110 166054 590730 201498
rect 590110 165818 590142 166054
rect 590378 165818 590462 166054
rect 590698 165818 590730 166054
rect 590110 165734 590730 165818
rect 590110 165498 590142 165734
rect 590378 165498 590462 165734
rect 590698 165498 590730 165734
rect 590110 130054 590730 165498
rect 590110 129818 590142 130054
rect 590378 129818 590462 130054
rect 590698 129818 590730 130054
rect 590110 129734 590730 129818
rect 590110 129498 590142 129734
rect 590378 129498 590462 129734
rect 590698 129498 590730 129734
rect 590110 94054 590730 129498
rect 590110 93818 590142 94054
rect 590378 93818 590462 94054
rect 590698 93818 590730 94054
rect 590110 93734 590730 93818
rect 590110 93498 590142 93734
rect 590378 93498 590462 93734
rect 590698 93498 590730 93734
rect 590110 58054 590730 93498
rect 590110 57818 590142 58054
rect 590378 57818 590462 58054
rect 590698 57818 590730 58054
rect 590110 57734 590730 57818
rect 590110 57498 590142 57734
rect 590378 57498 590462 57734
rect 590698 57498 590730 57734
rect 590110 22054 590730 57498
rect 590110 21818 590142 22054
rect 590378 21818 590462 22054
rect 590698 21818 590730 22054
rect 590110 21734 590730 21818
rect 590110 21498 590142 21734
rect 590378 21498 590462 21734
rect 590698 21498 590730 21734
rect 590110 -5146 590730 21498
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 673774 591690 710042
rect 591070 673538 591102 673774
rect 591338 673538 591422 673774
rect 591658 673538 591690 673774
rect 591070 673454 591690 673538
rect 591070 673218 591102 673454
rect 591338 673218 591422 673454
rect 591658 673218 591690 673454
rect 591070 637774 591690 673218
rect 591070 637538 591102 637774
rect 591338 637538 591422 637774
rect 591658 637538 591690 637774
rect 591070 637454 591690 637538
rect 591070 637218 591102 637454
rect 591338 637218 591422 637454
rect 591658 637218 591690 637454
rect 591070 601774 591690 637218
rect 591070 601538 591102 601774
rect 591338 601538 591422 601774
rect 591658 601538 591690 601774
rect 591070 601454 591690 601538
rect 591070 601218 591102 601454
rect 591338 601218 591422 601454
rect 591658 601218 591690 601454
rect 591070 565774 591690 601218
rect 591070 565538 591102 565774
rect 591338 565538 591422 565774
rect 591658 565538 591690 565774
rect 591070 565454 591690 565538
rect 591070 565218 591102 565454
rect 591338 565218 591422 565454
rect 591658 565218 591690 565454
rect 591070 529774 591690 565218
rect 591070 529538 591102 529774
rect 591338 529538 591422 529774
rect 591658 529538 591690 529774
rect 591070 529454 591690 529538
rect 591070 529218 591102 529454
rect 591338 529218 591422 529454
rect 591658 529218 591690 529454
rect 591070 493774 591690 529218
rect 591070 493538 591102 493774
rect 591338 493538 591422 493774
rect 591658 493538 591690 493774
rect 591070 493454 591690 493538
rect 591070 493218 591102 493454
rect 591338 493218 591422 493454
rect 591658 493218 591690 493454
rect 591070 457774 591690 493218
rect 591070 457538 591102 457774
rect 591338 457538 591422 457774
rect 591658 457538 591690 457774
rect 591070 457454 591690 457538
rect 591070 457218 591102 457454
rect 591338 457218 591422 457454
rect 591658 457218 591690 457454
rect 591070 421774 591690 457218
rect 591070 421538 591102 421774
rect 591338 421538 591422 421774
rect 591658 421538 591690 421774
rect 591070 421454 591690 421538
rect 591070 421218 591102 421454
rect 591338 421218 591422 421454
rect 591658 421218 591690 421454
rect 591070 385774 591690 421218
rect 591070 385538 591102 385774
rect 591338 385538 591422 385774
rect 591658 385538 591690 385774
rect 591070 385454 591690 385538
rect 591070 385218 591102 385454
rect 591338 385218 591422 385454
rect 591658 385218 591690 385454
rect 591070 349774 591690 385218
rect 591070 349538 591102 349774
rect 591338 349538 591422 349774
rect 591658 349538 591690 349774
rect 591070 349454 591690 349538
rect 591070 349218 591102 349454
rect 591338 349218 591422 349454
rect 591658 349218 591690 349454
rect 591070 313774 591690 349218
rect 591070 313538 591102 313774
rect 591338 313538 591422 313774
rect 591658 313538 591690 313774
rect 591070 313454 591690 313538
rect 591070 313218 591102 313454
rect 591338 313218 591422 313454
rect 591658 313218 591690 313454
rect 591070 277774 591690 313218
rect 591070 277538 591102 277774
rect 591338 277538 591422 277774
rect 591658 277538 591690 277774
rect 591070 277454 591690 277538
rect 591070 277218 591102 277454
rect 591338 277218 591422 277454
rect 591658 277218 591690 277454
rect 591070 241774 591690 277218
rect 591070 241538 591102 241774
rect 591338 241538 591422 241774
rect 591658 241538 591690 241774
rect 591070 241454 591690 241538
rect 591070 241218 591102 241454
rect 591338 241218 591422 241454
rect 591658 241218 591690 241454
rect 591070 205774 591690 241218
rect 591070 205538 591102 205774
rect 591338 205538 591422 205774
rect 591658 205538 591690 205774
rect 591070 205454 591690 205538
rect 591070 205218 591102 205454
rect 591338 205218 591422 205454
rect 591658 205218 591690 205454
rect 591070 169774 591690 205218
rect 591070 169538 591102 169774
rect 591338 169538 591422 169774
rect 591658 169538 591690 169774
rect 591070 169454 591690 169538
rect 591070 169218 591102 169454
rect 591338 169218 591422 169454
rect 591658 169218 591690 169454
rect 591070 133774 591690 169218
rect 591070 133538 591102 133774
rect 591338 133538 591422 133774
rect 591658 133538 591690 133774
rect 591070 133454 591690 133538
rect 591070 133218 591102 133454
rect 591338 133218 591422 133454
rect 591658 133218 591690 133454
rect 591070 97774 591690 133218
rect 591070 97538 591102 97774
rect 591338 97538 591422 97774
rect 591658 97538 591690 97774
rect 591070 97454 591690 97538
rect 591070 97218 591102 97454
rect 591338 97218 591422 97454
rect 591658 97218 591690 97454
rect 591070 61774 591690 97218
rect 591070 61538 591102 61774
rect 591338 61538 591422 61774
rect 591658 61538 591690 61774
rect 591070 61454 591690 61538
rect 591070 61218 591102 61454
rect 591338 61218 591422 61454
rect 591658 61218 591690 61454
rect 591070 25774 591690 61218
rect 591070 25538 591102 25774
rect 591338 25538 591422 25774
rect 591658 25538 591690 25774
rect 591070 25454 591690 25538
rect 591070 25218 591102 25454
rect 591338 25218 591422 25454
rect 591658 25218 591690 25454
rect 591070 -6106 591690 25218
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 677494 592650 711002
rect 592030 677258 592062 677494
rect 592298 677258 592382 677494
rect 592618 677258 592650 677494
rect 592030 677174 592650 677258
rect 592030 676938 592062 677174
rect 592298 676938 592382 677174
rect 592618 676938 592650 677174
rect 592030 641494 592650 676938
rect 592030 641258 592062 641494
rect 592298 641258 592382 641494
rect 592618 641258 592650 641494
rect 592030 641174 592650 641258
rect 592030 640938 592062 641174
rect 592298 640938 592382 641174
rect 592618 640938 592650 641174
rect 592030 605494 592650 640938
rect 592030 605258 592062 605494
rect 592298 605258 592382 605494
rect 592618 605258 592650 605494
rect 592030 605174 592650 605258
rect 592030 604938 592062 605174
rect 592298 604938 592382 605174
rect 592618 604938 592650 605174
rect 592030 569494 592650 604938
rect 592030 569258 592062 569494
rect 592298 569258 592382 569494
rect 592618 569258 592650 569494
rect 592030 569174 592650 569258
rect 592030 568938 592062 569174
rect 592298 568938 592382 569174
rect 592618 568938 592650 569174
rect 592030 533494 592650 568938
rect 592030 533258 592062 533494
rect 592298 533258 592382 533494
rect 592618 533258 592650 533494
rect 592030 533174 592650 533258
rect 592030 532938 592062 533174
rect 592298 532938 592382 533174
rect 592618 532938 592650 533174
rect 592030 497494 592650 532938
rect 592030 497258 592062 497494
rect 592298 497258 592382 497494
rect 592618 497258 592650 497494
rect 592030 497174 592650 497258
rect 592030 496938 592062 497174
rect 592298 496938 592382 497174
rect 592618 496938 592650 497174
rect 592030 461494 592650 496938
rect 592030 461258 592062 461494
rect 592298 461258 592382 461494
rect 592618 461258 592650 461494
rect 592030 461174 592650 461258
rect 592030 460938 592062 461174
rect 592298 460938 592382 461174
rect 592618 460938 592650 461174
rect 592030 425494 592650 460938
rect 592030 425258 592062 425494
rect 592298 425258 592382 425494
rect 592618 425258 592650 425494
rect 592030 425174 592650 425258
rect 592030 424938 592062 425174
rect 592298 424938 592382 425174
rect 592618 424938 592650 425174
rect 592030 389494 592650 424938
rect 592030 389258 592062 389494
rect 592298 389258 592382 389494
rect 592618 389258 592650 389494
rect 592030 389174 592650 389258
rect 592030 388938 592062 389174
rect 592298 388938 592382 389174
rect 592618 388938 592650 389174
rect 592030 353494 592650 388938
rect 592030 353258 592062 353494
rect 592298 353258 592382 353494
rect 592618 353258 592650 353494
rect 592030 353174 592650 353258
rect 592030 352938 592062 353174
rect 592298 352938 592382 353174
rect 592618 352938 592650 353174
rect 592030 317494 592650 352938
rect 592030 317258 592062 317494
rect 592298 317258 592382 317494
rect 592618 317258 592650 317494
rect 592030 317174 592650 317258
rect 592030 316938 592062 317174
rect 592298 316938 592382 317174
rect 592618 316938 592650 317174
rect 592030 281494 592650 316938
rect 592030 281258 592062 281494
rect 592298 281258 592382 281494
rect 592618 281258 592650 281494
rect 592030 281174 592650 281258
rect 592030 280938 592062 281174
rect 592298 280938 592382 281174
rect 592618 280938 592650 281174
rect 592030 245494 592650 280938
rect 592030 245258 592062 245494
rect 592298 245258 592382 245494
rect 592618 245258 592650 245494
rect 592030 245174 592650 245258
rect 592030 244938 592062 245174
rect 592298 244938 592382 245174
rect 592618 244938 592650 245174
rect 592030 209494 592650 244938
rect 592030 209258 592062 209494
rect 592298 209258 592382 209494
rect 592618 209258 592650 209494
rect 592030 209174 592650 209258
rect 592030 208938 592062 209174
rect 592298 208938 592382 209174
rect 592618 208938 592650 209174
rect 592030 173494 592650 208938
rect 592030 173258 592062 173494
rect 592298 173258 592382 173494
rect 592618 173258 592650 173494
rect 592030 173174 592650 173258
rect 592030 172938 592062 173174
rect 592298 172938 592382 173174
rect 592618 172938 592650 173174
rect 592030 137494 592650 172938
rect 592030 137258 592062 137494
rect 592298 137258 592382 137494
rect 592618 137258 592650 137494
rect 592030 137174 592650 137258
rect 592030 136938 592062 137174
rect 592298 136938 592382 137174
rect 592618 136938 592650 137174
rect 592030 101494 592650 136938
rect 592030 101258 592062 101494
rect 592298 101258 592382 101494
rect 592618 101258 592650 101494
rect 592030 101174 592650 101258
rect 592030 100938 592062 101174
rect 592298 100938 592382 101174
rect 592618 100938 592650 101174
rect 592030 65494 592650 100938
rect 592030 65258 592062 65494
rect 592298 65258 592382 65494
rect 592618 65258 592650 65494
rect 592030 65174 592650 65258
rect 592030 64938 592062 65174
rect 592298 64938 592382 65174
rect 592618 64938 592650 65174
rect 592030 29494 592650 64938
rect 592030 29258 592062 29494
rect 592298 29258 592382 29494
rect 592618 29258 592650 29494
rect 592030 29174 592650 29258
rect 592030 28938 592062 29174
rect 592298 28938 592382 29174
rect 592618 28938 592650 29174
rect 592030 -7066 592650 28938
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 677258 -8458 677494
rect -8374 677258 -8138 677494
rect -8694 676938 -8458 677174
rect -8374 676938 -8138 677174
rect -8694 641258 -8458 641494
rect -8374 641258 -8138 641494
rect -8694 640938 -8458 641174
rect -8374 640938 -8138 641174
rect -8694 605258 -8458 605494
rect -8374 605258 -8138 605494
rect -8694 604938 -8458 605174
rect -8374 604938 -8138 605174
rect -8694 569258 -8458 569494
rect -8374 569258 -8138 569494
rect -8694 568938 -8458 569174
rect -8374 568938 -8138 569174
rect -8694 533258 -8458 533494
rect -8374 533258 -8138 533494
rect -8694 532938 -8458 533174
rect -8374 532938 -8138 533174
rect -8694 497258 -8458 497494
rect -8374 497258 -8138 497494
rect -8694 496938 -8458 497174
rect -8374 496938 -8138 497174
rect -8694 461258 -8458 461494
rect -8374 461258 -8138 461494
rect -8694 460938 -8458 461174
rect -8374 460938 -8138 461174
rect -8694 425258 -8458 425494
rect -8374 425258 -8138 425494
rect -8694 424938 -8458 425174
rect -8374 424938 -8138 425174
rect -8694 389258 -8458 389494
rect -8374 389258 -8138 389494
rect -8694 388938 -8458 389174
rect -8374 388938 -8138 389174
rect -8694 353258 -8458 353494
rect -8374 353258 -8138 353494
rect -8694 352938 -8458 353174
rect -8374 352938 -8138 353174
rect -8694 317258 -8458 317494
rect -8374 317258 -8138 317494
rect -8694 316938 -8458 317174
rect -8374 316938 -8138 317174
rect -8694 281258 -8458 281494
rect -8374 281258 -8138 281494
rect -8694 280938 -8458 281174
rect -8374 280938 -8138 281174
rect -8694 245258 -8458 245494
rect -8374 245258 -8138 245494
rect -8694 244938 -8458 245174
rect -8374 244938 -8138 245174
rect -8694 209258 -8458 209494
rect -8374 209258 -8138 209494
rect -8694 208938 -8458 209174
rect -8374 208938 -8138 209174
rect -8694 173258 -8458 173494
rect -8374 173258 -8138 173494
rect -8694 172938 -8458 173174
rect -8374 172938 -8138 173174
rect -8694 137258 -8458 137494
rect -8374 137258 -8138 137494
rect -8694 136938 -8458 137174
rect -8374 136938 -8138 137174
rect -8694 101258 -8458 101494
rect -8374 101258 -8138 101494
rect -8694 100938 -8458 101174
rect -8374 100938 -8138 101174
rect -8694 65258 -8458 65494
rect -8374 65258 -8138 65494
rect -8694 64938 -8458 65174
rect -8374 64938 -8138 65174
rect -8694 29258 -8458 29494
rect -8374 29258 -8138 29494
rect -8694 28938 -8458 29174
rect -8374 28938 -8138 29174
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect -7734 673538 -7498 673774
rect -7414 673538 -7178 673774
rect -7734 673218 -7498 673454
rect -7414 673218 -7178 673454
rect -7734 637538 -7498 637774
rect -7414 637538 -7178 637774
rect -7734 637218 -7498 637454
rect -7414 637218 -7178 637454
rect -7734 601538 -7498 601774
rect -7414 601538 -7178 601774
rect -7734 601218 -7498 601454
rect -7414 601218 -7178 601454
rect -7734 565538 -7498 565774
rect -7414 565538 -7178 565774
rect -7734 565218 -7498 565454
rect -7414 565218 -7178 565454
rect -7734 529538 -7498 529774
rect -7414 529538 -7178 529774
rect -7734 529218 -7498 529454
rect -7414 529218 -7178 529454
rect -7734 493538 -7498 493774
rect -7414 493538 -7178 493774
rect -7734 493218 -7498 493454
rect -7414 493218 -7178 493454
rect -7734 457538 -7498 457774
rect -7414 457538 -7178 457774
rect -7734 457218 -7498 457454
rect -7414 457218 -7178 457454
rect -7734 421538 -7498 421774
rect -7414 421538 -7178 421774
rect -7734 421218 -7498 421454
rect -7414 421218 -7178 421454
rect -7734 385538 -7498 385774
rect -7414 385538 -7178 385774
rect -7734 385218 -7498 385454
rect -7414 385218 -7178 385454
rect -7734 349538 -7498 349774
rect -7414 349538 -7178 349774
rect -7734 349218 -7498 349454
rect -7414 349218 -7178 349454
rect -7734 313538 -7498 313774
rect -7414 313538 -7178 313774
rect -7734 313218 -7498 313454
rect -7414 313218 -7178 313454
rect -7734 277538 -7498 277774
rect -7414 277538 -7178 277774
rect -7734 277218 -7498 277454
rect -7414 277218 -7178 277454
rect -7734 241538 -7498 241774
rect -7414 241538 -7178 241774
rect -7734 241218 -7498 241454
rect -7414 241218 -7178 241454
rect -7734 205538 -7498 205774
rect -7414 205538 -7178 205774
rect -7734 205218 -7498 205454
rect -7414 205218 -7178 205454
rect -7734 169538 -7498 169774
rect -7414 169538 -7178 169774
rect -7734 169218 -7498 169454
rect -7414 169218 -7178 169454
rect -7734 133538 -7498 133774
rect -7414 133538 -7178 133774
rect -7734 133218 -7498 133454
rect -7414 133218 -7178 133454
rect -7734 97538 -7498 97774
rect -7414 97538 -7178 97774
rect -7734 97218 -7498 97454
rect -7414 97218 -7178 97454
rect -7734 61538 -7498 61774
rect -7414 61538 -7178 61774
rect -7734 61218 -7498 61454
rect -7414 61218 -7178 61454
rect -7734 25538 -7498 25774
rect -7414 25538 -7178 25774
rect -7734 25218 -7498 25454
rect -7414 25218 -7178 25454
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 669818 -6538 670054
rect -6454 669818 -6218 670054
rect -6774 669498 -6538 669734
rect -6454 669498 -6218 669734
rect -6774 633818 -6538 634054
rect -6454 633818 -6218 634054
rect -6774 633498 -6538 633734
rect -6454 633498 -6218 633734
rect -6774 597818 -6538 598054
rect -6454 597818 -6218 598054
rect -6774 597498 -6538 597734
rect -6454 597498 -6218 597734
rect -6774 561818 -6538 562054
rect -6454 561818 -6218 562054
rect -6774 561498 -6538 561734
rect -6454 561498 -6218 561734
rect -6774 525818 -6538 526054
rect -6454 525818 -6218 526054
rect -6774 525498 -6538 525734
rect -6454 525498 -6218 525734
rect -6774 489818 -6538 490054
rect -6454 489818 -6218 490054
rect -6774 489498 -6538 489734
rect -6454 489498 -6218 489734
rect -6774 453818 -6538 454054
rect -6454 453818 -6218 454054
rect -6774 453498 -6538 453734
rect -6454 453498 -6218 453734
rect -6774 417818 -6538 418054
rect -6454 417818 -6218 418054
rect -6774 417498 -6538 417734
rect -6454 417498 -6218 417734
rect -6774 381818 -6538 382054
rect -6454 381818 -6218 382054
rect -6774 381498 -6538 381734
rect -6454 381498 -6218 381734
rect -6774 345818 -6538 346054
rect -6454 345818 -6218 346054
rect -6774 345498 -6538 345734
rect -6454 345498 -6218 345734
rect -6774 309818 -6538 310054
rect -6454 309818 -6218 310054
rect -6774 309498 -6538 309734
rect -6454 309498 -6218 309734
rect -6774 273818 -6538 274054
rect -6454 273818 -6218 274054
rect -6774 273498 -6538 273734
rect -6454 273498 -6218 273734
rect -6774 237818 -6538 238054
rect -6454 237818 -6218 238054
rect -6774 237498 -6538 237734
rect -6454 237498 -6218 237734
rect -6774 201818 -6538 202054
rect -6454 201818 -6218 202054
rect -6774 201498 -6538 201734
rect -6454 201498 -6218 201734
rect -6774 165818 -6538 166054
rect -6454 165818 -6218 166054
rect -6774 165498 -6538 165734
rect -6454 165498 -6218 165734
rect -6774 129818 -6538 130054
rect -6454 129818 -6218 130054
rect -6774 129498 -6538 129734
rect -6454 129498 -6218 129734
rect -6774 93818 -6538 94054
rect -6454 93818 -6218 94054
rect -6774 93498 -6538 93734
rect -6454 93498 -6218 93734
rect -6774 57818 -6538 58054
rect -6454 57818 -6218 58054
rect -6774 57498 -6538 57734
rect -6454 57498 -6218 57734
rect -6774 21818 -6538 22054
rect -6454 21818 -6218 22054
rect -6774 21498 -6538 21734
rect -6454 21498 -6218 21734
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect -5814 666098 -5578 666334
rect -5494 666098 -5258 666334
rect -5814 665778 -5578 666014
rect -5494 665778 -5258 666014
rect -5814 630098 -5578 630334
rect -5494 630098 -5258 630334
rect -5814 629778 -5578 630014
rect -5494 629778 -5258 630014
rect -5814 594098 -5578 594334
rect -5494 594098 -5258 594334
rect -5814 593778 -5578 594014
rect -5494 593778 -5258 594014
rect -5814 558098 -5578 558334
rect -5494 558098 -5258 558334
rect -5814 557778 -5578 558014
rect -5494 557778 -5258 558014
rect -5814 522098 -5578 522334
rect -5494 522098 -5258 522334
rect -5814 521778 -5578 522014
rect -5494 521778 -5258 522014
rect -5814 486098 -5578 486334
rect -5494 486098 -5258 486334
rect -5814 485778 -5578 486014
rect -5494 485778 -5258 486014
rect -5814 450098 -5578 450334
rect -5494 450098 -5258 450334
rect -5814 449778 -5578 450014
rect -5494 449778 -5258 450014
rect -5814 414098 -5578 414334
rect -5494 414098 -5258 414334
rect -5814 413778 -5578 414014
rect -5494 413778 -5258 414014
rect -5814 378098 -5578 378334
rect -5494 378098 -5258 378334
rect -5814 377778 -5578 378014
rect -5494 377778 -5258 378014
rect -5814 342098 -5578 342334
rect -5494 342098 -5258 342334
rect -5814 341778 -5578 342014
rect -5494 341778 -5258 342014
rect -5814 306098 -5578 306334
rect -5494 306098 -5258 306334
rect -5814 305778 -5578 306014
rect -5494 305778 -5258 306014
rect -5814 270098 -5578 270334
rect -5494 270098 -5258 270334
rect -5814 269778 -5578 270014
rect -5494 269778 -5258 270014
rect -5814 234098 -5578 234334
rect -5494 234098 -5258 234334
rect -5814 233778 -5578 234014
rect -5494 233778 -5258 234014
rect -5814 198098 -5578 198334
rect -5494 198098 -5258 198334
rect -5814 197778 -5578 198014
rect -5494 197778 -5258 198014
rect -5814 162098 -5578 162334
rect -5494 162098 -5258 162334
rect -5814 161778 -5578 162014
rect -5494 161778 -5258 162014
rect -5814 126098 -5578 126334
rect -5494 126098 -5258 126334
rect -5814 125778 -5578 126014
rect -5494 125778 -5258 126014
rect -5814 90098 -5578 90334
rect -5494 90098 -5258 90334
rect -5814 89778 -5578 90014
rect -5494 89778 -5258 90014
rect -5814 54098 -5578 54334
rect -5494 54098 -5258 54334
rect -5814 53778 -5578 54014
rect -5494 53778 -5258 54014
rect -5814 18098 -5578 18334
rect -5494 18098 -5258 18334
rect -5814 17778 -5578 18014
rect -5494 17778 -5258 18014
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 698378 -4618 698614
rect -4534 698378 -4298 698614
rect -4854 698058 -4618 698294
rect -4534 698058 -4298 698294
rect -4854 662378 -4618 662614
rect -4534 662378 -4298 662614
rect -4854 662058 -4618 662294
rect -4534 662058 -4298 662294
rect -4854 626378 -4618 626614
rect -4534 626378 -4298 626614
rect -4854 626058 -4618 626294
rect -4534 626058 -4298 626294
rect -4854 590378 -4618 590614
rect -4534 590378 -4298 590614
rect -4854 590058 -4618 590294
rect -4534 590058 -4298 590294
rect -4854 554378 -4618 554614
rect -4534 554378 -4298 554614
rect -4854 554058 -4618 554294
rect -4534 554058 -4298 554294
rect -4854 518378 -4618 518614
rect -4534 518378 -4298 518614
rect -4854 518058 -4618 518294
rect -4534 518058 -4298 518294
rect -4854 482378 -4618 482614
rect -4534 482378 -4298 482614
rect -4854 482058 -4618 482294
rect -4534 482058 -4298 482294
rect -4854 446378 -4618 446614
rect -4534 446378 -4298 446614
rect -4854 446058 -4618 446294
rect -4534 446058 -4298 446294
rect -4854 410378 -4618 410614
rect -4534 410378 -4298 410614
rect -4854 410058 -4618 410294
rect -4534 410058 -4298 410294
rect -4854 374378 -4618 374614
rect -4534 374378 -4298 374614
rect -4854 374058 -4618 374294
rect -4534 374058 -4298 374294
rect -4854 338378 -4618 338614
rect -4534 338378 -4298 338614
rect -4854 338058 -4618 338294
rect -4534 338058 -4298 338294
rect -4854 302378 -4618 302614
rect -4534 302378 -4298 302614
rect -4854 302058 -4618 302294
rect -4534 302058 -4298 302294
rect -4854 266378 -4618 266614
rect -4534 266378 -4298 266614
rect -4854 266058 -4618 266294
rect -4534 266058 -4298 266294
rect -4854 230378 -4618 230614
rect -4534 230378 -4298 230614
rect -4854 230058 -4618 230294
rect -4534 230058 -4298 230294
rect -4854 194378 -4618 194614
rect -4534 194378 -4298 194614
rect -4854 194058 -4618 194294
rect -4534 194058 -4298 194294
rect -4854 158378 -4618 158614
rect -4534 158378 -4298 158614
rect -4854 158058 -4618 158294
rect -4534 158058 -4298 158294
rect -4854 122378 -4618 122614
rect -4534 122378 -4298 122614
rect -4854 122058 -4618 122294
rect -4534 122058 -4298 122294
rect -4854 86378 -4618 86614
rect -4534 86378 -4298 86614
rect -4854 86058 -4618 86294
rect -4534 86058 -4298 86294
rect -4854 50378 -4618 50614
rect -4534 50378 -4298 50614
rect -4854 50058 -4618 50294
rect -4534 50058 -4298 50294
rect -4854 14378 -4618 14614
rect -4534 14378 -4298 14614
rect -4854 14058 -4618 14294
rect -4534 14058 -4298 14294
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect -3894 694658 -3658 694894
rect -3574 694658 -3338 694894
rect -3894 694338 -3658 694574
rect -3574 694338 -3338 694574
rect -3894 658658 -3658 658894
rect -3574 658658 -3338 658894
rect -3894 658338 -3658 658574
rect -3574 658338 -3338 658574
rect -3894 622658 -3658 622894
rect -3574 622658 -3338 622894
rect -3894 622338 -3658 622574
rect -3574 622338 -3338 622574
rect -3894 586658 -3658 586894
rect -3574 586658 -3338 586894
rect -3894 586338 -3658 586574
rect -3574 586338 -3338 586574
rect -3894 550658 -3658 550894
rect -3574 550658 -3338 550894
rect -3894 550338 -3658 550574
rect -3574 550338 -3338 550574
rect -3894 514658 -3658 514894
rect -3574 514658 -3338 514894
rect -3894 514338 -3658 514574
rect -3574 514338 -3338 514574
rect -3894 478658 -3658 478894
rect -3574 478658 -3338 478894
rect -3894 478338 -3658 478574
rect -3574 478338 -3338 478574
rect -3894 442658 -3658 442894
rect -3574 442658 -3338 442894
rect -3894 442338 -3658 442574
rect -3574 442338 -3338 442574
rect -3894 406658 -3658 406894
rect -3574 406658 -3338 406894
rect -3894 406338 -3658 406574
rect -3574 406338 -3338 406574
rect -3894 370658 -3658 370894
rect -3574 370658 -3338 370894
rect -3894 370338 -3658 370574
rect -3574 370338 -3338 370574
rect -3894 334658 -3658 334894
rect -3574 334658 -3338 334894
rect -3894 334338 -3658 334574
rect -3574 334338 -3338 334574
rect -3894 298658 -3658 298894
rect -3574 298658 -3338 298894
rect -3894 298338 -3658 298574
rect -3574 298338 -3338 298574
rect -3894 262658 -3658 262894
rect -3574 262658 -3338 262894
rect -3894 262338 -3658 262574
rect -3574 262338 -3338 262574
rect -3894 226658 -3658 226894
rect -3574 226658 -3338 226894
rect -3894 226338 -3658 226574
rect -3574 226338 -3338 226574
rect -3894 190658 -3658 190894
rect -3574 190658 -3338 190894
rect -3894 190338 -3658 190574
rect -3574 190338 -3338 190574
rect -3894 154658 -3658 154894
rect -3574 154658 -3338 154894
rect -3894 154338 -3658 154574
rect -3574 154338 -3338 154574
rect -3894 118658 -3658 118894
rect -3574 118658 -3338 118894
rect -3894 118338 -3658 118574
rect -3574 118338 -3338 118574
rect -3894 82658 -3658 82894
rect -3574 82658 -3338 82894
rect -3894 82338 -3658 82574
rect -3574 82338 -3338 82574
rect -3894 46658 -3658 46894
rect -3574 46658 -3338 46894
rect -3894 46338 -3658 46574
rect -3574 46338 -3338 46574
rect -3894 10658 -3658 10894
rect -3574 10658 -3338 10894
rect -3894 10338 -3658 10574
rect -3574 10338 -3338 10574
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 690938 -2698 691174
rect -2614 690938 -2378 691174
rect -2934 690618 -2698 690854
rect -2614 690618 -2378 690854
rect -2934 654938 -2698 655174
rect -2614 654938 -2378 655174
rect -2934 654618 -2698 654854
rect -2614 654618 -2378 654854
rect -2934 618938 -2698 619174
rect -2614 618938 -2378 619174
rect -2934 618618 -2698 618854
rect -2614 618618 -2378 618854
rect -2934 582938 -2698 583174
rect -2614 582938 -2378 583174
rect -2934 582618 -2698 582854
rect -2614 582618 -2378 582854
rect -2934 546938 -2698 547174
rect -2614 546938 -2378 547174
rect -2934 546618 -2698 546854
rect -2614 546618 -2378 546854
rect -2934 510938 -2698 511174
rect -2614 510938 -2378 511174
rect -2934 510618 -2698 510854
rect -2614 510618 -2378 510854
rect -2934 474938 -2698 475174
rect -2614 474938 -2378 475174
rect -2934 474618 -2698 474854
rect -2614 474618 -2378 474854
rect -2934 438938 -2698 439174
rect -2614 438938 -2378 439174
rect -2934 438618 -2698 438854
rect -2614 438618 -2378 438854
rect -2934 402938 -2698 403174
rect -2614 402938 -2378 403174
rect -2934 402618 -2698 402854
rect -2614 402618 -2378 402854
rect -2934 366938 -2698 367174
rect -2614 366938 -2378 367174
rect -2934 366618 -2698 366854
rect -2614 366618 -2378 366854
rect -2934 330938 -2698 331174
rect -2614 330938 -2378 331174
rect -2934 330618 -2698 330854
rect -2614 330618 -2378 330854
rect -2934 294938 -2698 295174
rect -2614 294938 -2378 295174
rect -2934 294618 -2698 294854
rect -2614 294618 -2378 294854
rect -2934 258938 -2698 259174
rect -2614 258938 -2378 259174
rect -2934 258618 -2698 258854
rect -2614 258618 -2378 258854
rect -2934 222938 -2698 223174
rect -2614 222938 -2378 223174
rect -2934 222618 -2698 222854
rect -2614 222618 -2378 222854
rect -2934 186938 -2698 187174
rect -2614 186938 -2378 187174
rect -2934 186618 -2698 186854
rect -2614 186618 -2378 186854
rect -2934 150938 -2698 151174
rect -2614 150938 -2378 151174
rect -2934 150618 -2698 150854
rect -2614 150618 -2378 150854
rect -2934 114938 -2698 115174
rect -2614 114938 -2378 115174
rect -2934 114618 -2698 114854
rect -2614 114618 -2378 114854
rect -2934 78938 -2698 79174
rect -2614 78938 -2378 79174
rect -2934 78618 -2698 78854
rect -2614 78618 -2378 78854
rect -2934 42938 -2698 43174
rect -2614 42938 -2378 43174
rect -2934 42618 -2698 42854
rect -2614 42618 -2378 42854
rect -2934 6938 -2698 7174
rect -2614 6938 -2378 7174
rect -2934 6618 -2698 6854
rect -2614 6618 -2378 6854
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 5546 705562 5782 705798
rect 5866 705562 6102 705798
rect 5546 705242 5782 705478
rect 5866 705242 6102 705478
rect 5546 690938 5782 691174
rect 5866 690938 6102 691174
rect 5546 690618 5782 690854
rect 5866 690618 6102 690854
rect 5546 654938 5782 655174
rect 5866 654938 6102 655174
rect 5546 654618 5782 654854
rect 5866 654618 6102 654854
rect 5546 618938 5782 619174
rect 5866 618938 6102 619174
rect 5546 618618 5782 618854
rect 5866 618618 6102 618854
rect 5546 582938 5782 583174
rect 5866 582938 6102 583174
rect 5546 582618 5782 582854
rect 5866 582618 6102 582854
rect 5546 546938 5782 547174
rect 5866 546938 6102 547174
rect 5546 546618 5782 546854
rect 5866 546618 6102 546854
rect 5546 510938 5782 511174
rect 5866 510938 6102 511174
rect 5546 510618 5782 510854
rect 5866 510618 6102 510854
rect 5546 474938 5782 475174
rect 5866 474938 6102 475174
rect 5546 474618 5782 474854
rect 5866 474618 6102 474854
rect 5546 438938 5782 439174
rect 5866 438938 6102 439174
rect 5546 438618 5782 438854
rect 5866 438618 6102 438854
rect 5546 402938 5782 403174
rect 5866 402938 6102 403174
rect 5546 402618 5782 402854
rect 5866 402618 6102 402854
rect 5546 366938 5782 367174
rect 5866 366938 6102 367174
rect 5546 366618 5782 366854
rect 5866 366618 6102 366854
rect 5546 330938 5782 331174
rect 5866 330938 6102 331174
rect 5546 330618 5782 330854
rect 5866 330618 6102 330854
rect 5546 294938 5782 295174
rect 5866 294938 6102 295174
rect 5546 294618 5782 294854
rect 5866 294618 6102 294854
rect 5546 258938 5782 259174
rect 5866 258938 6102 259174
rect 5546 258618 5782 258854
rect 5866 258618 6102 258854
rect 5546 222938 5782 223174
rect 5866 222938 6102 223174
rect 5546 222618 5782 222854
rect 5866 222618 6102 222854
rect 5546 186938 5782 187174
rect 5866 186938 6102 187174
rect 5546 186618 5782 186854
rect 5866 186618 6102 186854
rect 5546 150938 5782 151174
rect 5866 150938 6102 151174
rect 5546 150618 5782 150854
rect 5866 150618 6102 150854
rect 5546 114938 5782 115174
rect 5866 114938 6102 115174
rect 5546 114618 5782 114854
rect 5866 114618 6102 114854
rect 5546 78938 5782 79174
rect 5866 78938 6102 79174
rect 5546 78618 5782 78854
rect 5866 78618 6102 78854
rect 5546 42938 5782 43174
rect 5866 42938 6102 43174
rect 5546 42618 5782 42854
rect 5866 42618 6102 42854
rect 5546 6938 5782 7174
rect 5866 6938 6102 7174
rect 5546 6618 5782 6854
rect 5866 6618 6102 6854
rect 5546 -1542 5782 -1306
rect 5866 -1542 6102 -1306
rect 5546 -1862 5782 -1626
rect 5866 -1862 6102 -1626
rect 9266 706522 9502 706758
rect 9586 706522 9822 706758
rect 9266 706202 9502 706438
rect 9586 706202 9822 706438
rect 9266 694658 9502 694894
rect 9586 694658 9822 694894
rect 9266 694338 9502 694574
rect 9586 694338 9822 694574
rect 12986 707482 13222 707718
rect 13306 707482 13542 707718
rect 12986 707162 13222 707398
rect 13306 707162 13542 707398
rect 12986 698378 13222 698614
rect 13306 698378 13542 698614
rect 12986 698058 13222 698294
rect 13306 698058 13542 698294
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 41546 705562 41782 705798
rect 41866 705562 42102 705798
rect 41546 705242 41782 705478
rect 41866 705242 42102 705478
rect 41546 690938 41782 691174
rect 41866 690938 42102 691174
rect 41546 690618 41782 690854
rect 41866 690618 42102 690854
rect 45266 706522 45502 706758
rect 45586 706522 45822 706758
rect 45266 706202 45502 706438
rect 45586 706202 45822 706438
rect 45266 694658 45502 694894
rect 45586 694658 45822 694894
rect 45266 694338 45502 694574
rect 45586 694338 45822 694574
rect 48986 707482 49222 707718
rect 49306 707482 49542 707718
rect 48986 707162 49222 707398
rect 49306 707162 49542 707398
rect 48986 698378 49222 698614
rect 49306 698378 49542 698614
rect 48986 698058 49222 698294
rect 49306 698058 49542 698294
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 77546 705562 77782 705798
rect 77866 705562 78102 705798
rect 77546 705242 77782 705478
rect 77866 705242 78102 705478
rect 77546 690938 77782 691174
rect 77866 690938 78102 691174
rect 77546 690618 77782 690854
rect 77866 690618 78102 690854
rect 81266 706522 81502 706758
rect 81586 706522 81822 706758
rect 81266 706202 81502 706438
rect 81586 706202 81822 706438
rect 81266 694658 81502 694894
rect 81586 694658 81822 694894
rect 81266 694338 81502 694574
rect 81586 694338 81822 694574
rect 84986 707482 85222 707718
rect 85306 707482 85542 707718
rect 84986 707162 85222 707398
rect 85306 707162 85542 707398
rect 84986 698378 85222 698614
rect 85306 698378 85542 698614
rect 84986 698058 85222 698294
rect 85306 698058 85542 698294
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 113546 705562 113782 705798
rect 113866 705562 114102 705798
rect 113546 705242 113782 705478
rect 113866 705242 114102 705478
rect 113546 690938 113782 691174
rect 113866 690938 114102 691174
rect 113546 690618 113782 690854
rect 113866 690618 114102 690854
rect 117266 706522 117502 706758
rect 117586 706522 117822 706758
rect 117266 706202 117502 706438
rect 117586 706202 117822 706438
rect 117266 694658 117502 694894
rect 117586 694658 117822 694894
rect 117266 694338 117502 694574
rect 117586 694338 117822 694574
rect 120986 707482 121222 707718
rect 121306 707482 121542 707718
rect 120986 707162 121222 707398
rect 121306 707162 121542 707398
rect 120986 698378 121222 698614
rect 121306 698378 121542 698614
rect 120986 698058 121222 698294
rect 121306 698058 121542 698294
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 149546 705562 149782 705798
rect 149866 705562 150102 705798
rect 149546 705242 149782 705478
rect 149866 705242 150102 705478
rect 149546 690938 149782 691174
rect 149866 690938 150102 691174
rect 149546 690618 149782 690854
rect 149866 690618 150102 690854
rect 153266 706522 153502 706758
rect 153586 706522 153822 706758
rect 153266 706202 153502 706438
rect 153586 706202 153822 706438
rect 153266 694658 153502 694894
rect 153586 694658 153822 694894
rect 153266 694338 153502 694574
rect 153586 694338 153822 694574
rect 156986 707482 157222 707718
rect 157306 707482 157542 707718
rect 156986 707162 157222 707398
rect 157306 707162 157542 707398
rect 156986 698378 157222 698614
rect 157306 698378 157542 698614
rect 156986 698058 157222 698294
rect 157306 698058 157542 698294
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 185546 705562 185782 705798
rect 185866 705562 186102 705798
rect 185546 705242 185782 705478
rect 185866 705242 186102 705478
rect 185546 690938 185782 691174
rect 185866 690938 186102 691174
rect 185546 690618 185782 690854
rect 185866 690618 186102 690854
rect 189266 706522 189502 706758
rect 189586 706522 189822 706758
rect 189266 706202 189502 706438
rect 189586 706202 189822 706438
rect 189266 694658 189502 694894
rect 189586 694658 189822 694894
rect 189266 694338 189502 694574
rect 189586 694338 189822 694574
rect 192986 707482 193222 707718
rect 193306 707482 193542 707718
rect 192986 707162 193222 707398
rect 193306 707162 193542 707398
rect 192986 698378 193222 698614
rect 193306 698378 193542 698614
rect 192986 698058 193222 698294
rect 193306 698058 193542 698294
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 221546 705562 221782 705798
rect 221866 705562 222102 705798
rect 221546 705242 221782 705478
rect 221866 705242 222102 705478
rect 221546 690938 221782 691174
rect 221866 690938 222102 691174
rect 221546 690618 221782 690854
rect 221866 690618 222102 690854
rect 225266 706522 225502 706758
rect 225586 706522 225822 706758
rect 225266 706202 225502 706438
rect 225586 706202 225822 706438
rect 225266 694658 225502 694894
rect 225586 694658 225822 694894
rect 225266 694338 225502 694574
rect 225586 694338 225822 694574
rect 228986 707482 229222 707718
rect 229306 707482 229542 707718
rect 228986 707162 229222 707398
rect 229306 707162 229542 707398
rect 228986 698378 229222 698614
rect 229306 698378 229542 698614
rect 228986 698058 229222 698294
rect 229306 698058 229542 698294
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 257546 705562 257782 705798
rect 257866 705562 258102 705798
rect 257546 705242 257782 705478
rect 257866 705242 258102 705478
rect 257546 690938 257782 691174
rect 257866 690938 258102 691174
rect 257546 690618 257782 690854
rect 257866 690618 258102 690854
rect 261266 706522 261502 706758
rect 261586 706522 261822 706758
rect 261266 706202 261502 706438
rect 261586 706202 261822 706438
rect 261266 694658 261502 694894
rect 261586 694658 261822 694894
rect 261266 694338 261502 694574
rect 261586 694338 261822 694574
rect 264986 707482 265222 707718
rect 265306 707482 265542 707718
rect 264986 707162 265222 707398
rect 265306 707162 265542 707398
rect 264986 698378 265222 698614
rect 265306 698378 265542 698614
rect 264986 698058 265222 698294
rect 265306 698058 265542 698294
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 293546 705562 293782 705798
rect 293866 705562 294102 705798
rect 293546 705242 293782 705478
rect 293866 705242 294102 705478
rect 293546 690938 293782 691174
rect 293866 690938 294102 691174
rect 293546 690618 293782 690854
rect 293866 690618 294102 690854
rect 297266 706522 297502 706758
rect 297586 706522 297822 706758
rect 297266 706202 297502 706438
rect 297586 706202 297822 706438
rect 297266 694658 297502 694894
rect 297586 694658 297822 694894
rect 297266 694338 297502 694574
rect 297586 694338 297822 694574
rect 300986 707482 301222 707718
rect 301306 707482 301542 707718
rect 300986 707162 301222 707398
rect 301306 707162 301542 707398
rect 300986 698378 301222 698614
rect 301306 698378 301542 698614
rect 300986 698058 301222 698294
rect 301306 698058 301542 698294
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 329546 705562 329782 705798
rect 329866 705562 330102 705798
rect 329546 705242 329782 705478
rect 329866 705242 330102 705478
rect 329546 690938 329782 691174
rect 329866 690938 330102 691174
rect 329546 690618 329782 690854
rect 329866 690618 330102 690854
rect 333266 706522 333502 706758
rect 333586 706522 333822 706758
rect 333266 706202 333502 706438
rect 333586 706202 333822 706438
rect 333266 694658 333502 694894
rect 333586 694658 333822 694894
rect 333266 694338 333502 694574
rect 333586 694338 333822 694574
rect 336986 707482 337222 707718
rect 337306 707482 337542 707718
rect 336986 707162 337222 707398
rect 337306 707162 337542 707398
rect 336986 698378 337222 698614
rect 337306 698378 337542 698614
rect 336986 698058 337222 698294
rect 337306 698058 337542 698294
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 365546 705562 365782 705798
rect 365866 705562 366102 705798
rect 365546 705242 365782 705478
rect 365866 705242 366102 705478
rect 365546 690938 365782 691174
rect 365866 690938 366102 691174
rect 365546 690618 365782 690854
rect 365866 690618 366102 690854
rect 369266 706522 369502 706758
rect 369586 706522 369822 706758
rect 369266 706202 369502 706438
rect 369586 706202 369822 706438
rect 369266 694658 369502 694894
rect 369586 694658 369822 694894
rect 369266 694338 369502 694574
rect 369586 694338 369822 694574
rect 372986 707482 373222 707718
rect 373306 707482 373542 707718
rect 372986 707162 373222 707398
rect 373306 707162 373542 707398
rect 372986 698378 373222 698614
rect 373306 698378 373542 698614
rect 372986 698058 373222 698294
rect 373306 698058 373542 698294
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 401546 705562 401782 705798
rect 401866 705562 402102 705798
rect 401546 705242 401782 705478
rect 401866 705242 402102 705478
rect 401546 690938 401782 691174
rect 401866 690938 402102 691174
rect 401546 690618 401782 690854
rect 401866 690618 402102 690854
rect 405266 706522 405502 706758
rect 405586 706522 405822 706758
rect 405266 706202 405502 706438
rect 405586 706202 405822 706438
rect 405266 694658 405502 694894
rect 405586 694658 405822 694894
rect 405266 694338 405502 694574
rect 405586 694338 405822 694574
rect 408986 707482 409222 707718
rect 409306 707482 409542 707718
rect 408986 707162 409222 707398
rect 409306 707162 409542 707398
rect 408986 698378 409222 698614
rect 409306 698378 409542 698614
rect 408986 698058 409222 698294
rect 409306 698058 409542 698294
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 437546 705562 437782 705798
rect 437866 705562 438102 705798
rect 437546 705242 437782 705478
rect 437866 705242 438102 705478
rect 437546 690938 437782 691174
rect 437866 690938 438102 691174
rect 437546 690618 437782 690854
rect 437866 690618 438102 690854
rect 441266 706522 441502 706758
rect 441586 706522 441822 706758
rect 441266 706202 441502 706438
rect 441586 706202 441822 706438
rect 441266 694658 441502 694894
rect 441586 694658 441822 694894
rect 441266 694338 441502 694574
rect 441586 694338 441822 694574
rect 444986 707482 445222 707718
rect 445306 707482 445542 707718
rect 444986 707162 445222 707398
rect 445306 707162 445542 707398
rect 444986 698378 445222 698614
rect 445306 698378 445542 698614
rect 444986 698058 445222 698294
rect 445306 698058 445542 698294
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 473546 705562 473782 705798
rect 473866 705562 474102 705798
rect 473546 705242 473782 705478
rect 473866 705242 474102 705478
rect 473546 690938 473782 691174
rect 473866 690938 474102 691174
rect 473546 690618 473782 690854
rect 473866 690618 474102 690854
rect 477266 706522 477502 706758
rect 477586 706522 477822 706758
rect 477266 706202 477502 706438
rect 477586 706202 477822 706438
rect 477266 694658 477502 694894
rect 477586 694658 477822 694894
rect 477266 694338 477502 694574
rect 477586 694338 477822 694574
rect 480986 707482 481222 707718
rect 481306 707482 481542 707718
rect 480986 707162 481222 707398
rect 481306 707162 481542 707398
rect 480986 698378 481222 698614
rect 481306 698378 481542 698614
rect 480986 698058 481222 698294
rect 481306 698058 481542 698294
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 509546 705562 509782 705798
rect 509866 705562 510102 705798
rect 509546 705242 509782 705478
rect 509866 705242 510102 705478
rect 509546 690938 509782 691174
rect 509866 690938 510102 691174
rect 509546 690618 509782 690854
rect 509866 690618 510102 690854
rect 513266 706522 513502 706758
rect 513586 706522 513822 706758
rect 513266 706202 513502 706438
rect 513586 706202 513822 706438
rect 513266 694658 513502 694894
rect 513586 694658 513822 694894
rect 513266 694338 513502 694574
rect 513586 694338 513822 694574
rect 516986 707482 517222 707718
rect 517306 707482 517542 707718
rect 516986 707162 517222 707398
rect 517306 707162 517542 707398
rect 516986 698378 517222 698614
rect 517306 698378 517542 698614
rect 516986 698058 517222 698294
rect 517306 698058 517542 698294
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 545546 705562 545782 705798
rect 545866 705562 546102 705798
rect 545546 705242 545782 705478
rect 545866 705242 546102 705478
rect 545546 690938 545782 691174
rect 545866 690938 546102 691174
rect 545546 690618 545782 690854
rect 545866 690618 546102 690854
rect 549266 706522 549502 706758
rect 549586 706522 549822 706758
rect 549266 706202 549502 706438
rect 549586 706202 549822 706438
rect 549266 694658 549502 694894
rect 549586 694658 549822 694894
rect 549266 694338 549502 694574
rect 549586 694338 549822 694574
rect 552986 707482 553222 707718
rect 553306 707482 553542 707718
rect 552986 707162 553222 707398
rect 553306 707162 553542 707398
rect 552986 698378 553222 698614
rect 553306 698378 553542 698614
rect 552986 698058 553222 698294
rect 553306 698058 553542 698294
rect 567866 711322 568102 711558
rect 568186 711322 568422 711558
rect 567866 711002 568102 711238
rect 568186 711002 568422 711238
rect 9266 658658 9502 658894
rect 9586 658658 9822 658894
rect 9266 658338 9502 658574
rect 9586 658338 9822 658574
rect 567866 677258 568102 677494
rect 568186 677258 568422 677494
rect 567866 676938 568102 677174
rect 568186 676938 568422 677174
rect 31610 654938 31846 655174
rect 31610 654618 31846 654854
rect 62330 654938 62566 655174
rect 62330 654618 62566 654854
rect 93050 654938 93286 655174
rect 93050 654618 93286 654854
rect 123770 654938 124006 655174
rect 123770 654618 124006 654854
rect 154490 654938 154726 655174
rect 154490 654618 154726 654854
rect 185210 654938 185446 655174
rect 185210 654618 185446 654854
rect 215930 654938 216166 655174
rect 215930 654618 216166 654854
rect 246650 654938 246886 655174
rect 246650 654618 246886 654854
rect 277370 654938 277606 655174
rect 277370 654618 277606 654854
rect 308090 654938 308326 655174
rect 308090 654618 308326 654854
rect 338810 654938 339046 655174
rect 338810 654618 339046 654854
rect 369530 654938 369766 655174
rect 369530 654618 369766 654854
rect 400250 654938 400486 655174
rect 400250 654618 400486 654854
rect 430970 654938 431206 655174
rect 430970 654618 431206 654854
rect 461690 654938 461926 655174
rect 461690 654618 461926 654854
rect 492410 654938 492646 655174
rect 492410 654618 492646 654854
rect 523130 654938 523366 655174
rect 523130 654618 523366 654854
rect 553850 654938 554086 655174
rect 553850 654618 554086 654854
rect 16250 651218 16486 651454
rect 16250 650898 16486 651134
rect 46970 651218 47206 651454
rect 46970 650898 47206 651134
rect 77690 651218 77926 651454
rect 77690 650898 77926 651134
rect 108410 651218 108646 651454
rect 108410 650898 108646 651134
rect 139130 651218 139366 651454
rect 139130 650898 139366 651134
rect 169850 651218 170086 651454
rect 169850 650898 170086 651134
rect 200570 651218 200806 651454
rect 200570 650898 200806 651134
rect 231290 651218 231526 651454
rect 231290 650898 231526 651134
rect 262010 651218 262246 651454
rect 262010 650898 262246 651134
rect 292730 651218 292966 651454
rect 292730 650898 292966 651134
rect 323450 651218 323686 651454
rect 323450 650898 323686 651134
rect 354170 651218 354406 651454
rect 354170 650898 354406 651134
rect 384890 651218 385126 651454
rect 384890 650898 385126 651134
rect 415610 651218 415846 651454
rect 415610 650898 415846 651134
rect 446330 651218 446566 651454
rect 446330 650898 446566 651134
rect 477050 651218 477286 651454
rect 477050 650898 477286 651134
rect 507770 651218 508006 651454
rect 507770 650898 508006 651134
rect 538490 651218 538726 651454
rect 538490 650898 538726 651134
rect 9266 622658 9502 622894
rect 9586 622658 9822 622894
rect 9266 622338 9502 622574
rect 9586 622338 9822 622574
rect 567866 641258 568102 641494
rect 568186 641258 568422 641494
rect 567866 640938 568102 641174
rect 568186 640938 568422 641174
rect 31610 618938 31846 619174
rect 31610 618618 31846 618854
rect 62330 618938 62566 619174
rect 62330 618618 62566 618854
rect 93050 618938 93286 619174
rect 93050 618618 93286 618854
rect 123770 618938 124006 619174
rect 123770 618618 124006 618854
rect 154490 618938 154726 619174
rect 154490 618618 154726 618854
rect 185210 618938 185446 619174
rect 185210 618618 185446 618854
rect 215930 618938 216166 619174
rect 215930 618618 216166 618854
rect 246650 618938 246886 619174
rect 246650 618618 246886 618854
rect 277370 618938 277606 619174
rect 277370 618618 277606 618854
rect 308090 618938 308326 619174
rect 308090 618618 308326 618854
rect 338810 618938 339046 619174
rect 338810 618618 339046 618854
rect 369530 618938 369766 619174
rect 369530 618618 369766 618854
rect 400250 618938 400486 619174
rect 400250 618618 400486 618854
rect 430970 618938 431206 619174
rect 430970 618618 431206 618854
rect 461690 618938 461926 619174
rect 461690 618618 461926 618854
rect 492410 618938 492646 619174
rect 492410 618618 492646 618854
rect 523130 618938 523366 619174
rect 523130 618618 523366 618854
rect 553850 618938 554086 619174
rect 553850 618618 554086 618854
rect 16250 615218 16486 615454
rect 16250 614898 16486 615134
rect 46970 615218 47206 615454
rect 46970 614898 47206 615134
rect 77690 615218 77926 615454
rect 77690 614898 77926 615134
rect 108410 615218 108646 615454
rect 108410 614898 108646 615134
rect 139130 615218 139366 615454
rect 139130 614898 139366 615134
rect 169850 615218 170086 615454
rect 169850 614898 170086 615134
rect 200570 615218 200806 615454
rect 200570 614898 200806 615134
rect 231290 615218 231526 615454
rect 231290 614898 231526 615134
rect 262010 615218 262246 615454
rect 262010 614898 262246 615134
rect 292730 615218 292966 615454
rect 292730 614898 292966 615134
rect 323450 615218 323686 615454
rect 323450 614898 323686 615134
rect 354170 615218 354406 615454
rect 354170 614898 354406 615134
rect 384890 615218 385126 615454
rect 384890 614898 385126 615134
rect 415610 615218 415846 615454
rect 415610 614898 415846 615134
rect 446330 615218 446566 615454
rect 446330 614898 446566 615134
rect 477050 615218 477286 615454
rect 477050 614898 477286 615134
rect 507770 615218 508006 615454
rect 507770 614898 508006 615134
rect 538490 615218 538726 615454
rect 538490 614898 538726 615134
rect 9266 586658 9502 586894
rect 9586 586658 9822 586894
rect 9266 586338 9502 586574
rect 9586 586338 9822 586574
rect 567866 605258 568102 605494
rect 568186 605258 568422 605494
rect 567866 604938 568102 605174
rect 568186 604938 568422 605174
rect 31610 582938 31846 583174
rect 31610 582618 31846 582854
rect 62330 582938 62566 583174
rect 62330 582618 62566 582854
rect 93050 582938 93286 583174
rect 93050 582618 93286 582854
rect 123770 582938 124006 583174
rect 123770 582618 124006 582854
rect 154490 582938 154726 583174
rect 154490 582618 154726 582854
rect 185210 582938 185446 583174
rect 185210 582618 185446 582854
rect 215930 582938 216166 583174
rect 215930 582618 216166 582854
rect 246650 582938 246886 583174
rect 246650 582618 246886 582854
rect 277370 582938 277606 583174
rect 277370 582618 277606 582854
rect 308090 582938 308326 583174
rect 308090 582618 308326 582854
rect 338810 582938 339046 583174
rect 338810 582618 339046 582854
rect 369530 582938 369766 583174
rect 369530 582618 369766 582854
rect 400250 582938 400486 583174
rect 400250 582618 400486 582854
rect 430970 582938 431206 583174
rect 430970 582618 431206 582854
rect 461690 582938 461926 583174
rect 461690 582618 461926 582854
rect 492410 582938 492646 583174
rect 492410 582618 492646 582854
rect 523130 582938 523366 583174
rect 523130 582618 523366 582854
rect 553850 582938 554086 583174
rect 553850 582618 554086 582854
rect 16250 579218 16486 579454
rect 16250 578898 16486 579134
rect 46970 579218 47206 579454
rect 46970 578898 47206 579134
rect 77690 579218 77926 579454
rect 77690 578898 77926 579134
rect 108410 579218 108646 579454
rect 108410 578898 108646 579134
rect 139130 579218 139366 579454
rect 139130 578898 139366 579134
rect 169850 579218 170086 579454
rect 169850 578898 170086 579134
rect 200570 579218 200806 579454
rect 200570 578898 200806 579134
rect 231290 579218 231526 579454
rect 231290 578898 231526 579134
rect 262010 579218 262246 579454
rect 262010 578898 262246 579134
rect 292730 579218 292966 579454
rect 292730 578898 292966 579134
rect 323450 579218 323686 579454
rect 323450 578898 323686 579134
rect 354170 579218 354406 579454
rect 354170 578898 354406 579134
rect 384890 579218 385126 579454
rect 384890 578898 385126 579134
rect 415610 579218 415846 579454
rect 415610 578898 415846 579134
rect 446330 579218 446566 579454
rect 446330 578898 446566 579134
rect 477050 579218 477286 579454
rect 477050 578898 477286 579134
rect 507770 579218 508006 579454
rect 507770 578898 508006 579134
rect 538490 579218 538726 579454
rect 538490 578898 538726 579134
rect 9266 550658 9502 550894
rect 9586 550658 9822 550894
rect 9266 550338 9502 550574
rect 9586 550338 9822 550574
rect 567866 569258 568102 569494
rect 568186 569258 568422 569494
rect 567866 568938 568102 569174
rect 568186 568938 568422 569174
rect 31610 546938 31846 547174
rect 31610 546618 31846 546854
rect 62330 546938 62566 547174
rect 62330 546618 62566 546854
rect 93050 546938 93286 547174
rect 93050 546618 93286 546854
rect 123770 546938 124006 547174
rect 123770 546618 124006 546854
rect 154490 546938 154726 547174
rect 154490 546618 154726 546854
rect 185210 546938 185446 547174
rect 185210 546618 185446 546854
rect 215930 546938 216166 547174
rect 215930 546618 216166 546854
rect 246650 546938 246886 547174
rect 246650 546618 246886 546854
rect 277370 546938 277606 547174
rect 277370 546618 277606 546854
rect 308090 546938 308326 547174
rect 308090 546618 308326 546854
rect 338810 546938 339046 547174
rect 338810 546618 339046 546854
rect 369530 546938 369766 547174
rect 369530 546618 369766 546854
rect 400250 546938 400486 547174
rect 400250 546618 400486 546854
rect 430970 546938 431206 547174
rect 430970 546618 431206 546854
rect 461690 546938 461926 547174
rect 461690 546618 461926 546854
rect 492410 546938 492646 547174
rect 492410 546618 492646 546854
rect 523130 546938 523366 547174
rect 523130 546618 523366 546854
rect 553850 546938 554086 547174
rect 553850 546618 554086 546854
rect 16250 543218 16486 543454
rect 16250 542898 16486 543134
rect 46970 543218 47206 543454
rect 46970 542898 47206 543134
rect 77690 543218 77926 543454
rect 77690 542898 77926 543134
rect 108410 543218 108646 543454
rect 108410 542898 108646 543134
rect 139130 543218 139366 543454
rect 139130 542898 139366 543134
rect 169850 543218 170086 543454
rect 169850 542898 170086 543134
rect 200570 543218 200806 543454
rect 200570 542898 200806 543134
rect 231290 543218 231526 543454
rect 231290 542898 231526 543134
rect 262010 543218 262246 543454
rect 262010 542898 262246 543134
rect 292730 543218 292966 543454
rect 292730 542898 292966 543134
rect 323450 543218 323686 543454
rect 323450 542898 323686 543134
rect 354170 543218 354406 543454
rect 354170 542898 354406 543134
rect 384890 543218 385126 543454
rect 384890 542898 385126 543134
rect 415610 543218 415846 543454
rect 415610 542898 415846 543134
rect 446330 543218 446566 543454
rect 446330 542898 446566 543134
rect 477050 543218 477286 543454
rect 477050 542898 477286 543134
rect 507770 543218 508006 543454
rect 507770 542898 508006 543134
rect 538490 543218 538726 543454
rect 538490 542898 538726 543134
rect 9266 514658 9502 514894
rect 9586 514658 9822 514894
rect 9266 514338 9502 514574
rect 9586 514338 9822 514574
rect 567866 533258 568102 533494
rect 568186 533258 568422 533494
rect 567866 532938 568102 533174
rect 568186 532938 568422 533174
rect 31610 510938 31846 511174
rect 31610 510618 31846 510854
rect 62330 510938 62566 511174
rect 62330 510618 62566 510854
rect 93050 510938 93286 511174
rect 93050 510618 93286 510854
rect 123770 510938 124006 511174
rect 123770 510618 124006 510854
rect 154490 510938 154726 511174
rect 154490 510618 154726 510854
rect 185210 510938 185446 511174
rect 185210 510618 185446 510854
rect 215930 510938 216166 511174
rect 215930 510618 216166 510854
rect 246650 510938 246886 511174
rect 246650 510618 246886 510854
rect 277370 510938 277606 511174
rect 277370 510618 277606 510854
rect 308090 510938 308326 511174
rect 308090 510618 308326 510854
rect 338810 510938 339046 511174
rect 338810 510618 339046 510854
rect 369530 510938 369766 511174
rect 369530 510618 369766 510854
rect 400250 510938 400486 511174
rect 400250 510618 400486 510854
rect 430970 510938 431206 511174
rect 430970 510618 431206 510854
rect 461690 510938 461926 511174
rect 461690 510618 461926 510854
rect 492410 510938 492646 511174
rect 492410 510618 492646 510854
rect 523130 510938 523366 511174
rect 523130 510618 523366 510854
rect 553850 510938 554086 511174
rect 553850 510618 554086 510854
rect 16250 507218 16486 507454
rect 16250 506898 16486 507134
rect 46970 507218 47206 507454
rect 46970 506898 47206 507134
rect 77690 507218 77926 507454
rect 77690 506898 77926 507134
rect 108410 507218 108646 507454
rect 108410 506898 108646 507134
rect 139130 507218 139366 507454
rect 139130 506898 139366 507134
rect 169850 507218 170086 507454
rect 169850 506898 170086 507134
rect 200570 507218 200806 507454
rect 200570 506898 200806 507134
rect 231290 507218 231526 507454
rect 231290 506898 231526 507134
rect 262010 507218 262246 507454
rect 262010 506898 262246 507134
rect 292730 507218 292966 507454
rect 292730 506898 292966 507134
rect 323450 507218 323686 507454
rect 323450 506898 323686 507134
rect 354170 507218 354406 507454
rect 354170 506898 354406 507134
rect 384890 507218 385126 507454
rect 384890 506898 385126 507134
rect 415610 507218 415846 507454
rect 415610 506898 415846 507134
rect 446330 507218 446566 507454
rect 446330 506898 446566 507134
rect 477050 507218 477286 507454
rect 477050 506898 477286 507134
rect 507770 507218 508006 507454
rect 507770 506898 508006 507134
rect 538490 507218 538726 507454
rect 538490 506898 538726 507134
rect 9266 478658 9502 478894
rect 9586 478658 9822 478894
rect 9266 478338 9502 478574
rect 9586 478338 9822 478574
rect 567866 497258 568102 497494
rect 568186 497258 568422 497494
rect 567866 496938 568102 497174
rect 568186 496938 568422 497174
rect 31610 474938 31846 475174
rect 31610 474618 31846 474854
rect 62330 474938 62566 475174
rect 62330 474618 62566 474854
rect 93050 474938 93286 475174
rect 93050 474618 93286 474854
rect 123770 474938 124006 475174
rect 123770 474618 124006 474854
rect 154490 474938 154726 475174
rect 154490 474618 154726 474854
rect 185210 474938 185446 475174
rect 185210 474618 185446 474854
rect 215930 474938 216166 475174
rect 215930 474618 216166 474854
rect 246650 474938 246886 475174
rect 246650 474618 246886 474854
rect 277370 474938 277606 475174
rect 277370 474618 277606 474854
rect 308090 474938 308326 475174
rect 308090 474618 308326 474854
rect 338810 474938 339046 475174
rect 338810 474618 339046 474854
rect 369530 474938 369766 475174
rect 369530 474618 369766 474854
rect 400250 474938 400486 475174
rect 400250 474618 400486 474854
rect 430970 474938 431206 475174
rect 430970 474618 431206 474854
rect 461690 474938 461926 475174
rect 461690 474618 461926 474854
rect 492410 474938 492646 475174
rect 492410 474618 492646 474854
rect 523130 474938 523366 475174
rect 523130 474618 523366 474854
rect 553850 474938 554086 475174
rect 553850 474618 554086 474854
rect 16250 471218 16486 471454
rect 16250 470898 16486 471134
rect 46970 471218 47206 471454
rect 46970 470898 47206 471134
rect 77690 471218 77926 471454
rect 77690 470898 77926 471134
rect 108410 471218 108646 471454
rect 108410 470898 108646 471134
rect 139130 471218 139366 471454
rect 139130 470898 139366 471134
rect 169850 471218 170086 471454
rect 169850 470898 170086 471134
rect 200570 471218 200806 471454
rect 200570 470898 200806 471134
rect 231290 471218 231526 471454
rect 231290 470898 231526 471134
rect 262010 471218 262246 471454
rect 262010 470898 262246 471134
rect 292730 471218 292966 471454
rect 292730 470898 292966 471134
rect 323450 471218 323686 471454
rect 323450 470898 323686 471134
rect 354170 471218 354406 471454
rect 354170 470898 354406 471134
rect 384890 471218 385126 471454
rect 384890 470898 385126 471134
rect 415610 471218 415846 471454
rect 415610 470898 415846 471134
rect 446330 471218 446566 471454
rect 446330 470898 446566 471134
rect 477050 471218 477286 471454
rect 477050 470898 477286 471134
rect 507770 471218 508006 471454
rect 507770 470898 508006 471134
rect 538490 471218 538726 471454
rect 538490 470898 538726 471134
rect 9266 442658 9502 442894
rect 9586 442658 9822 442894
rect 9266 442338 9502 442574
rect 9586 442338 9822 442574
rect 567866 461258 568102 461494
rect 568186 461258 568422 461494
rect 567866 460938 568102 461174
rect 568186 460938 568422 461174
rect 31610 438938 31846 439174
rect 31610 438618 31846 438854
rect 62330 438938 62566 439174
rect 62330 438618 62566 438854
rect 93050 438938 93286 439174
rect 93050 438618 93286 438854
rect 123770 438938 124006 439174
rect 123770 438618 124006 438854
rect 154490 438938 154726 439174
rect 154490 438618 154726 438854
rect 185210 438938 185446 439174
rect 185210 438618 185446 438854
rect 215930 438938 216166 439174
rect 215930 438618 216166 438854
rect 246650 438938 246886 439174
rect 246650 438618 246886 438854
rect 277370 438938 277606 439174
rect 277370 438618 277606 438854
rect 308090 438938 308326 439174
rect 308090 438618 308326 438854
rect 338810 438938 339046 439174
rect 338810 438618 339046 438854
rect 369530 438938 369766 439174
rect 369530 438618 369766 438854
rect 400250 438938 400486 439174
rect 400250 438618 400486 438854
rect 430970 438938 431206 439174
rect 430970 438618 431206 438854
rect 461690 438938 461926 439174
rect 461690 438618 461926 438854
rect 492410 438938 492646 439174
rect 492410 438618 492646 438854
rect 523130 438938 523366 439174
rect 523130 438618 523366 438854
rect 553850 438938 554086 439174
rect 553850 438618 554086 438854
rect 16250 435218 16486 435454
rect 16250 434898 16486 435134
rect 46970 435218 47206 435454
rect 46970 434898 47206 435134
rect 77690 435218 77926 435454
rect 77690 434898 77926 435134
rect 108410 435218 108646 435454
rect 108410 434898 108646 435134
rect 139130 435218 139366 435454
rect 139130 434898 139366 435134
rect 169850 435218 170086 435454
rect 169850 434898 170086 435134
rect 200570 435218 200806 435454
rect 200570 434898 200806 435134
rect 231290 435218 231526 435454
rect 231290 434898 231526 435134
rect 262010 435218 262246 435454
rect 262010 434898 262246 435134
rect 292730 435218 292966 435454
rect 292730 434898 292966 435134
rect 323450 435218 323686 435454
rect 323450 434898 323686 435134
rect 354170 435218 354406 435454
rect 354170 434898 354406 435134
rect 384890 435218 385126 435454
rect 384890 434898 385126 435134
rect 415610 435218 415846 435454
rect 415610 434898 415846 435134
rect 446330 435218 446566 435454
rect 446330 434898 446566 435134
rect 477050 435218 477286 435454
rect 477050 434898 477286 435134
rect 507770 435218 508006 435454
rect 507770 434898 508006 435134
rect 538490 435218 538726 435454
rect 538490 434898 538726 435134
rect 9266 406658 9502 406894
rect 9586 406658 9822 406894
rect 9266 406338 9502 406574
rect 9586 406338 9822 406574
rect 567866 425258 568102 425494
rect 568186 425258 568422 425494
rect 567866 424938 568102 425174
rect 568186 424938 568422 425174
rect 31610 402938 31846 403174
rect 31610 402618 31846 402854
rect 62330 402938 62566 403174
rect 62330 402618 62566 402854
rect 93050 402938 93286 403174
rect 93050 402618 93286 402854
rect 123770 402938 124006 403174
rect 123770 402618 124006 402854
rect 154490 402938 154726 403174
rect 154490 402618 154726 402854
rect 185210 402938 185446 403174
rect 185210 402618 185446 402854
rect 215930 402938 216166 403174
rect 215930 402618 216166 402854
rect 246650 402938 246886 403174
rect 246650 402618 246886 402854
rect 277370 402938 277606 403174
rect 277370 402618 277606 402854
rect 308090 402938 308326 403174
rect 308090 402618 308326 402854
rect 338810 402938 339046 403174
rect 338810 402618 339046 402854
rect 369530 402938 369766 403174
rect 369530 402618 369766 402854
rect 400250 402938 400486 403174
rect 400250 402618 400486 402854
rect 430970 402938 431206 403174
rect 430970 402618 431206 402854
rect 461690 402938 461926 403174
rect 461690 402618 461926 402854
rect 492410 402938 492646 403174
rect 492410 402618 492646 402854
rect 523130 402938 523366 403174
rect 523130 402618 523366 402854
rect 553850 402938 554086 403174
rect 553850 402618 554086 402854
rect 16250 399218 16486 399454
rect 16250 398898 16486 399134
rect 46970 399218 47206 399454
rect 46970 398898 47206 399134
rect 77690 399218 77926 399454
rect 77690 398898 77926 399134
rect 108410 399218 108646 399454
rect 108410 398898 108646 399134
rect 139130 399218 139366 399454
rect 139130 398898 139366 399134
rect 169850 399218 170086 399454
rect 169850 398898 170086 399134
rect 200570 399218 200806 399454
rect 200570 398898 200806 399134
rect 231290 399218 231526 399454
rect 231290 398898 231526 399134
rect 262010 399218 262246 399454
rect 262010 398898 262246 399134
rect 292730 399218 292966 399454
rect 292730 398898 292966 399134
rect 323450 399218 323686 399454
rect 323450 398898 323686 399134
rect 354170 399218 354406 399454
rect 354170 398898 354406 399134
rect 384890 399218 385126 399454
rect 384890 398898 385126 399134
rect 415610 399218 415846 399454
rect 415610 398898 415846 399134
rect 446330 399218 446566 399454
rect 446330 398898 446566 399134
rect 477050 399218 477286 399454
rect 477050 398898 477286 399134
rect 507770 399218 508006 399454
rect 507770 398898 508006 399134
rect 538490 399218 538726 399454
rect 538490 398898 538726 399134
rect 9266 370658 9502 370894
rect 9586 370658 9822 370894
rect 9266 370338 9502 370574
rect 9586 370338 9822 370574
rect 567866 389258 568102 389494
rect 568186 389258 568422 389494
rect 567866 388938 568102 389174
rect 568186 388938 568422 389174
rect 31610 366938 31846 367174
rect 31610 366618 31846 366854
rect 62330 366938 62566 367174
rect 62330 366618 62566 366854
rect 93050 366938 93286 367174
rect 93050 366618 93286 366854
rect 123770 366938 124006 367174
rect 123770 366618 124006 366854
rect 154490 366938 154726 367174
rect 154490 366618 154726 366854
rect 185210 366938 185446 367174
rect 185210 366618 185446 366854
rect 215930 366938 216166 367174
rect 215930 366618 216166 366854
rect 246650 366938 246886 367174
rect 246650 366618 246886 366854
rect 277370 366938 277606 367174
rect 277370 366618 277606 366854
rect 308090 366938 308326 367174
rect 308090 366618 308326 366854
rect 338810 366938 339046 367174
rect 338810 366618 339046 366854
rect 369530 366938 369766 367174
rect 369530 366618 369766 366854
rect 400250 366938 400486 367174
rect 400250 366618 400486 366854
rect 430970 366938 431206 367174
rect 430970 366618 431206 366854
rect 461690 366938 461926 367174
rect 461690 366618 461926 366854
rect 492410 366938 492646 367174
rect 492410 366618 492646 366854
rect 523130 366938 523366 367174
rect 523130 366618 523366 366854
rect 553850 366938 554086 367174
rect 553850 366618 554086 366854
rect 16250 363218 16486 363454
rect 16250 362898 16486 363134
rect 46970 363218 47206 363454
rect 46970 362898 47206 363134
rect 77690 363218 77926 363454
rect 77690 362898 77926 363134
rect 108410 363218 108646 363454
rect 108410 362898 108646 363134
rect 139130 363218 139366 363454
rect 139130 362898 139366 363134
rect 169850 363218 170086 363454
rect 169850 362898 170086 363134
rect 200570 363218 200806 363454
rect 200570 362898 200806 363134
rect 231290 363218 231526 363454
rect 231290 362898 231526 363134
rect 262010 363218 262246 363454
rect 262010 362898 262246 363134
rect 292730 363218 292966 363454
rect 292730 362898 292966 363134
rect 323450 363218 323686 363454
rect 323450 362898 323686 363134
rect 354170 363218 354406 363454
rect 354170 362898 354406 363134
rect 384890 363218 385126 363454
rect 384890 362898 385126 363134
rect 415610 363218 415846 363454
rect 415610 362898 415846 363134
rect 446330 363218 446566 363454
rect 446330 362898 446566 363134
rect 477050 363218 477286 363454
rect 477050 362898 477286 363134
rect 507770 363218 508006 363454
rect 507770 362898 508006 363134
rect 538490 363218 538726 363454
rect 538490 362898 538726 363134
rect 9266 334658 9502 334894
rect 9586 334658 9822 334894
rect 9266 334338 9502 334574
rect 9586 334338 9822 334574
rect 567866 353258 568102 353494
rect 568186 353258 568422 353494
rect 567866 352938 568102 353174
rect 568186 352938 568422 353174
rect 31610 330938 31846 331174
rect 31610 330618 31846 330854
rect 62330 330938 62566 331174
rect 62330 330618 62566 330854
rect 93050 330938 93286 331174
rect 93050 330618 93286 330854
rect 123770 330938 124006 331174
rect 123770 330618 124006 330854
rect 154490 330938 154726 331174
rect 154490 330618 154726 330854
rect 185210 330938 185446 331174
rect 185210 330618 185446 330854
rect 215930 330938 216166 331174
rect 215930 330618 216166 330854
rect 246650 330938 246886 331174
rect 246650 330618 246886 330854
rect 277370 330938 277606 331174
rect 277370 330618 277606 330854
rect 308090 330938 308326 331174
rect 308090 330618 308326 330854
rect 338810 330938 339046 331174
rect 338810 330618 339046 330854
rect 369530 330938 369766 331174
rect 369530 330618 369766 330854
rect 400250 330938 400486 331174
rect 400250 330618 400486 330854
rect 430970 330938 431206 331174
rect 430970 330618 431206 330854
rect 461690 330938 461926 331174
rect 461690 330618 461926 330854
rect 492410 330938 492646 331174
rect 492410 330618 492646 330854
rect 523130 330938 523366 331174
rect 523130 330618 523366 330854
rect 553850 330938 554086 331174
rect 553850 330618 554086 330854
rect 16250 327218 16486 327454
rect 16250 326898 16486 327134
rect 46970 327218 47206 327454
rect 46970 326898 47206 327134
rect 77690 327218 77926 327454
rect 77690 326898 77926 327134
rect 108410 327218 108646 327454
rect 108410 326898 108646 327134
rect 139130 327218 139366 327454
rect 139130 326898 139366 327134
rect 169850 327218 170086 327454
rect 169850 326898 170086 327134
rect 200570 327218 200806 327454
rect 200570 326898 200806 327134
rect 231290 327218 231526 327454
rect 231290 326898 231526 327134
rect 262010 327218 262246 327454
rect 262010 326898 262246 327134
rect 292730 327218 292966 327454
rect 292730 326898 292966 327134
rect 323450 327218 323686 327454
rect 323450 326898 323686 327134
rect 354170 327218 354406 327454
rect 354170 326898 354406 327134
rect 384890 327218 385126 327454
rect 384890 326898 385126 327134
rect 415610 327218 415846 327454
rect 415610 326898 415846 327134
rect 446330 327218 446566 327454
rect 446330 326898 446566 327134
rect 477050 327218 477286 327454
rect 477050 326898 477286 327134
rect 507770 327218 508006 327454
rect 507770 326898 508006 327134
rect 538490 327218 538726 327454
rect 538490 326898 538726 327134
rect 9266 298658 9502 298894
rect 9586 298658 9822 298894
rect 9266 298338 9502 298574
rect 9586 298338 9822 298574
rect 567866 317258 568102 317494
rect 568186 317258 568422 317494
rect 567866 316938 568102 317174
rect 568186 316938 568422 317174
rect 31610 294938 31846 295174
rect 31610 294618 31846 294854
rect 62330 294938 62566 295174
rect 62330 294618 62566 294854
rect 93050 294938 93286 295174
rect 93050 294618 93286 294854
rect 123770 294938 124006 295174
rect 123770 294618 124006 294854
rect 154490 294938 154726 295174
rect 154490 294618 154726 294854
rect 185210 294938 185446 295174
rect 185210 294618 185446 294854
rect 215930 294938 216166 295174
rect 215930 294618 216166 294854
rect 246650 294938 246886 295174
rect 246650 294618 246886 294854
rect 277370 294938 277606 295174
rect 277370 294618 277606 294854
rect 308090 294938 308326 295174
rect 308090 294618 308326 294854
rect 338810 294938 339046 295174
rect 338810 294618 339046 294854
rect 369530 294938 369766 295174
rect 369530 294618 369766 294854
rect 400250 294938 400486 295174
rect 400250 294618 400486 294854
rect 430970 294938 431206 295174
rect 430970 294618 431206 294854
rect 461690 294938 461926 295174
rect 461690 294618 461926 294854
rect 492410 294938 492646 295174
rect 492410 294618 492646 294854
rect 523130 294938 523366 295174
rect 523130 294618 523366 294854
rect 553850 294938 554086 295174
rect 553850 294618 554086 294854
rect 16250 291218 16486 291454
rect 16250 290898 16486 291134
rect 46970 291218 47206 291454
rect 46970 290898 47206 291134
rect 77690 291218 77926 291454
rect 77690 290898 77926 291134
rect 108410 291218 108646 291454
rect 108410 290898 108646 291134
rect 139130 291218 139366 291454
rect 139130 290898 139366 291134
rect 169850 291218 170086 291454
rect 169850 290898 170086 291134
rect 200570 291218 200806 291454
rect 200570 290898 200806 291134
rect 231290 291218 231526 291454
rect 231290 290898 231526 291134
rect 262010 291218 262246 291454
rect 262010 290898 262246 291134
rect 292730 291218 292966 291454
rect 292730 290898 292966 291134
rect 323450 291218 323686 291454
rect 323450 290898 323686 291134
rect 354170 291218 354406 291454
rect 354170 290898 354406 291134
rect 384890 291218 385126 291454
rect 384890 290898 385126 291134
rect 415610 291218 415846 291454
rect 415610 290898 415846 291134
rect 446330 291218 446566 291454
rect 446330 290898 446566 291134
rect 477050 291218 477286 291454
rect 477050 290898 477286 291134
rect 507770 291218 508006 291454
rect 507770 290898 508006 291134
rect 538490 291218 538726 291454
rect 538490 290898 538726 291134
rect 9266 262658 9502 262894
rect 9586 262658 9822 262894
rect 9266 262338 9502 262574
rect 9586 262338 9822 262574
rect 567866 281258 568102 281494
rect 568186 281258 568422 281494
rect 567866 280938 568102 281174
rect 568186 280938 568422 281174
rect 31610 258938 31846 259174
rect 31610 258618 31846 258854
rect 62330 258938 62566 259174
rect 62330 258618 62566 258854
rect 93050 258938 93286 259174
rect 93050 258618 93286 258854
rect 123770 258938 124006 259174
rect 123770 258618 124006 258854
rect 154490 258938 154726 259174
rect 154490 258618 154726 258854
rect 185210 258938 185446 259174
rect 185210 258618 185446 258854
rect 215930 258938 216166 259174
rect 215930 258618 216166 258854
rect 246650 258938 246886 259174
rect 246650 258618 246886 258854
rect 277370 258938 277606 259174
rect 277370 258618 277606 258854
rect 308090 258938 308326 259174
rect 308090 258618 308326 258854
rect 338810 258938 339046 259174
rect 338810 258618 339046 258854
rect 369530 258938 369766 259174
rect 369530 258618 369766 258854
rect 400250 258938 400486 259174
rect 400250 258618 400486 258854
rect 430970 258938 431206 259174
rect 430970 258618 431206 258854
rect 461690 258938 461926 259174
rect 461690 258618 461926 258854
rect 492410 258938 492646 259174
rect 492410 258618 492646 258854
rect 523130 258938 523366 259174
rect 523130 258618 523366 258854
rect 553850 258938 554086 259174
rect 553850 258618 554086 258854
rect 16250 255218 16486 255454
rect 16250 254898 16486 255134
rect 46970 255218 47206 255454
rect 46970 254898 47206 255134
rect 77690 255218 77926 255454
rect 77690 254898 77926 255134
rect 108410 255218 108646 255454
rect 108410 254898 108646 255134
rect 139130 255218 139366 255454
rect 139130 254898 139366 255134
rect 169850 255218 170086 255454
rect 169850 254898 170086 255134
rect 200570 255218 200806 255454
rect 200570 254898 200806 255134
rect 231290 255218 231526 255454
rect 231290 254898 231526 255134
rect 262010 255218 262246 255454
rect 262010 254898 262246 255134
rect 292730 255218 292966 255454
rect 292730 254898 292966 255134
rect 323450 255218 323686 255454
rect 323450 254898 323686 255134
rect 354170 255218 354406 255454
rect 354170 254898 354406 255134
rect 384890 255218 385126 255454
rect 384890 254898 385126 255134
rect 415610 255218 415846 255454
rect 415610 254898 415846 255134
rect 446330 255218 446566 255454
rect 446330 254898 446566 255134
rect 477050 255218 477286 255454
rect 477050 254898 477286 255134
rect 507770 255218 508006 255454
rect 507770 254898 508006 255134
rect 538490 255218 538726 255454
rect 538490 254898 538726 255134
rect 9266 226658 9502 226894
rect 9586 226658 9822 226894
rect 9266 226338 9502 226574
rect 9586 226338 9822 226574
rect 567866 245258 568102 245494
rect 568186 245258 568422 245494
rect 567866 244938 568102 245174
rect 568186 244938 568422 245174
rect 31610 222938 31846 223174
rect 31610 222618 31846 222854
rect 62330 222938 62566 223174
rect 62330 222618 62566 222854
rect 93050 222938 93286 223174
rect 93050 222618 93286 222854
rect 123770 222938 124006 223174
rect 123770 222618 124006 222854
rect 154490 222938 154726 223174
rect 154490 222618 154726 222854
rect 185210 222938 185446 223174
rect 185210 222618 185446 222854
rect 215930 222938 216166 223174
rect 215930 222618 216166 222854
rect 246650 222938 246886 223174
rect 246650 222618 246886 222854
rect 277370 222938 277606 223174
rect 277370 222618 277606 222854
rect 308090 222938 308326 223174
rect 308090 222618 308326 222854
rect 338810 222938 339046 223174
rect 338810 222618 339046 222854
rect 369530 222938 369766 223174
rect 369530 222618 369766 222854
rect 400250 222938 400486 223174
rect 400250 222618 400486 222854
rect 430970 222938 431206 223174
rect 430970 222618 431206 222854
rect 461690 222938 461926 223174
rect 461690 222618 461926 222854
rect 492410 222938 492646 223174
rect 492410 222618 492646 222854
rect 523130 222938 523366 223174
rect 523130 222618 523366 222854
rect 553850 222938 554086 223174
rect 553850 222618 554086 222854
rect 16250 219218 16486 219454
rect 16250 218898 16486 219134
rect 46970 219218 47206 219454
rect 46970 218898 47206 219134
rect 77690 219218 77926 219454
rect 77690 218898 77926 219134
rect 108410 219218 108646 219454
rect 108410 218898 108646 219134
rect 139130 219218 139366 219454
rect 139130 218898 139366 219134
rect 169850 219218 170086 219454
rect 169850 218898 170086 219134
rect 200570 219218 200806 219454
rect 200570 218898 200806 219134
rect 231290 219218 231526 219454
rect 231290 218898 231526 219134
rect 262010 219218 262246 219454
rect 262010 218898 262246 219134
rect 292730 219218 292966 219454
rect 292730 218898 292966 219134
rect 323450 219218 323686 219454
rect 323450 218898 323686 219134
rect 354170 219218 354406 219454
rect 354170 218898 354406 219134
rect 384890 219218 385126 219454
rect 384890 218898 385126 219134
rect 415610 219218 415846 219454
rect 415610 218898 415846 219134
rect 446330 219218 446566 219454
rect 446330 218898 446566 219134
rect 477050 219218 477286 219454
rect 477050 218898 477286 219134
rect 507770 219218 508006 219454
rect 507770 218898 508006 219134
rect 538490 219218 538726 219454
rect 538490 218898 538726 219134
rect 9266 190658 9502 190894
rect 9586 190658 9822 190894
rect 9266 190338 9502 190574
rect 9586 190338 9822 190574
rect 567866 209258 568102 209494
rect 568186 209258 568422 209494
rect 567866 208938 568102 209174
rect 568186 208938 568422 209174
rect 31610 186938 31846 187174
rect 31610 186618 31846 186854
rect 62330 186938 62566 187174
rect 62330 186618 62566 186854
rect 93050 186938 93286 187174
rect 93050 186618 93286 186854
rect 123770 186938 124006 187174
rect 123770 186618 124006 186854
rect 154490 186938 154726 187174
rect 154490 186618 154726 186854
rect 185210 186938 185446 187174
rect 185210 186618 185446 186854
rect 215930 186938 216166 187174
rect 215930 186618 216166 186854
rect 246650 186938 246886 187174
rect 246650 186618 246886 186854
rect 277370 186938 277606 187174
rect 277370 186618 277606 186854
rect 308090 186938 308326 187174
rect 308090 186618 308326 186854
rect 338810 186938 339046 187174
rect 338810 186618 339046 186854
rect 369530 186938 369766 187174
rect 369530 186618 369766 186854
rect 400250 186938 400486 187174
rect 400250 186618 400486 186854
rect 430970 186938 431206 187174
rect 430970 186618 431206 186854
rect 461690 186938 461926 187174
rect 461690 186618 461926 186854
rect 492410 186938 492646 187174
rect 492410 186618 492646 186854
rect 523130 186938 523366 187174
rect 523130 186618 523366 186854
rect 553850 186938 554086 187174
rect 553850 186618 554086 186854
rect 16250 183218 16486 183454
rect 16250 182898 16486 183134
rect 46970 183218 47206 183454
rect 46970 182898 47206 183134
rect 77690 183218 77926 183454
rect 77690 182898 77926 183134
rect 108410 183218 108646 183454
rect 108410 182898 108646 183134
rect 139130 183218 139366 183454
rect 139130 182898 139366 183134
rect 169850 183218 170086 183454
rect 169850 182898 170086 183134
rect 200570 183218 200806 183454
rect 200570 182898 200806 183134
rect 231290 183218 231526 183454
rect 231290 182898 231526 183134
rect 262010 183218 262246 183454
rect 262010 182898 262246 183134
rect 292730 183218 292966 183454
rect 292730 182898 292966 183134
rect 323450 183218 323686 183454
rect 323450 182898 323686 183134
rect 354170 183218 354406 183454
rect 354170 182898 354406 183134
rect 384890 183218 385126 183454
rect 384890 182898 385126 183134
rect 415610 183218 415846 183454
rect 415610 182898 415846 183134
rect 446330 183218 446566 183454
rect 446330 182898 446566 183134
rect 477050 183218 477286 183454
rect 477050 182898 477286 183134
rect 507770 183218 508006 183454
rect 507770 182898 508006 183134
rect 538490 183218 538726 183454
rect 538490 182898 538726 183134
rect 9266 154658 9502 154894
rect 9586 154658 9822 154894
rect 9266 154338 9502 154574
rect 9586 154338 9822 154574
rect 567866 173258 568102 173494
rect 568186 173258 568422 173494
rect 567866 172938 568102 173174
rect 568186 172938 568422 173174
rect 31610 150938 31846 151174
rect 31610 150618 31846 150854
rect 62330 150938 62566 151174
rect 62330 150618 62566 150854
rect 93050 150938 93286 151174
rect 93050 150618 93286 150854
rect 123770 150938 124006 151174
rect 123770 150618 124006 150854
rect 154490 150938 154726 151174
rect 154490 150618 154726 150854
rect 185210 150938 185446 151174
rect 185210 150618 185446 150854
rect 215930 150938 216166 151174
rect 215930 150618 216166 150854
rect 246650 150938 246886 151174
rect 246650 150618 246886 150854
rect 277370 150938 277606 151174
rect 277370 150618 277606 150854
rect 308090 150938 308326 151174
rect 308090 150618 308326 150854
rect 338810 150938 339046 151174
rect 338810 150618 339046 150854
rect 369530 150938 369766 151174
rect 369530 150618 369766 150854
rect 400250 150938 400486 151174
rect 400250 150618 400486 150854
rect 430970 150938 431206 151174
rect 430970 150618 431206 150854
rect 461690 150938 461926 151174
rect 461690 150618 461926 150854
rect 492410 150938 492646 151174
rect 492410 150618 492646 150854
rect 523130 150938 523366 151174
rect 523130 150618 523366 150854
rect 553850 150938 554086 151174
rect 553850 150618 554086 150854
rect 16250 147218 16486 147454
rect 16250 146898 16486 147134
rect 46970 147218 47206 147454
rect 46970 146898 47206 147134
rect 77690 147218 77926 147454
rect 77690 146898 77926 147134
rect 108410 147218 108646 147454
rect 108410 146898 108646 147134
rect 139130 147218 139366 147454
rect 139130 146898 139366 147134
rect 169850 147218 170086 147454
rect 169850 146898 170086 147134
rect 200570 147218 200806 147454
rect 200570 146898 200806 147134
rect 231290 147218 231526 147454
rect 231290 146898 231526 147134
rect 262010 147218 262246 147454
rect 262010 146898 262246 147134
rect 292730 147218 292966 147454
rect 292730 146898 292966 147134
rect 323450 147218 323686 147454
rect 323450 146898 323686 147134
rect 354170 147218 354406 147454
rect 354170 146898 354406 147134
rect 384890 147218 385126 147454
rect 384890 146898 385126 147134
rect 415610 147218 415846 147454
rect 415610 146898 415846 147134
rect 446330 147218 446566 147454
rect 446330 146898 446566 147134
rect 477050 147218 477286 147454
rect 477050 146898 477286 147134
rect 507770 147218 508006 147454
rect 507770 146898 508006 147134
rect 538490 147218 538726 147454
rect 538490 146898 538726 147134
rect 9266 118658 9502 118894
rect 9586 118658 9822 118894
rect 9266 118338 9502 118574
rect 9586 118338 9822 118574
rect 567866 137258 568102 137494
rect 568186 137258 568422 137494
rect 567866 136938 568102 137174
rect 568186 136938 568422 137174
rect 31610 114938 31846 115174
rect 31610 114618 31846 114854
rect 62330 114938 62566 115174
rect 62330 114618 62566 114854
rect 93050 114938 93286 115174
rect 93050 114618 93286 114854
rect 123770 114938 124006 115174
rect 123770 114618 124006 114854
rect 154490 114938 154726 115174
rect 154490 114618 154726 114854
rect 185210 114938 185446 115174
rect 185210 114618 185446 114854
rect 215930 114938 216166 115174
rect 215930 114618 216166 114854
rect 246650 114938 246886 115174
rect 246650 114618 246886 114854
rect 277370 114938 277606 115174
rect 277370 114618 277606 114854
rect 308090 114938 308326 115174
rect 308090 114618 308326 114854
rect 338810 114938 339046 115174
rect 338810 114618 339046 114854
rect 369530 114938 369766 115174
rect 369530 114618 369766 114854
rect 400250 114938 400486 115174
rect 400250 114618 400486 114854
rect 430970 114938 431206 115174
rect 430970 114618 431206 114854
rect 461690 114938 461926 115174
rect 461690 114618 461926 114854
rect 492410 114938 492646 115174
rect 492410 114618 492646 114854
rect 523130 114938 523366 115174
rect 523130 114618 523366 114854
rect 553850 114938 554086 115174
rect 553850 114618 554086 114854
rect 16250 111218 16486 111454
rect 16250 110898 16486 111134
rect 46970 111218 47206 111454
rect 46970 110898 47206 111134
rect 77690 111218 77926 111454
rect 77690 110898 77926 111134
rect 108410 111218 108646 111454
rect 108410 110898 108646 111134
rect 139130 111218 139366 111454
rect 139130 110898 139366 111134
rect 169850 111218 170086 111454
rect 169850 110898 170086 111134
rect 200570 111218 200806 111454
rect 200570 110898 200806 111134
rect 231290 111218 231526 111454
rect 231290 110898 231526 111134
rect 262010 111218 262246 111454
rect 262010 110898 262246 111134
rect 292730 111218 292966 111454
rect 292730 110898 292966 111134
rect 323450 111218 323686 111454
rect 323450 110898 323686 111134
rect 354170 111218 354406 111454
rect 354170 110898 354406 111134
rect 384890 111218 385126 111454
rect 384890 110898 385126 111134
rect 415610 111218 415846 111454
rect 415610 110898 415846 111134
rect 446330 111218 446566 111454
rect 446330 110898 446566 111134
rect 477050 111218 477286 111454
rect 477050 110898 477286 111134
rect 507770 111218 508006 111454
rect 507770 110898 508006 111134
rect 538490 111218 538726 111454
rect 538490 110898 538726 111134
rect 9266 82658 9502 82894
rect 9586 82658 9822 82894
rect 9266 82338 9502 82574
rect 9586 82338 9822 82574
rect 567866 101258 568102 101494
rect 568186 101258 568422 101494
rect 567866 100938 568102 101174
rect 568186 100938 568422 101174
rect 31610 78938 31846 79174
rect 31610 78618 31846 78854
rect 62330 78938 62566 79174
rect 62330 78618 62566 78854
rect 93050 78938 93286 79174
rect 93050 78618 93286 78854
rect 123770 78938 124006 79174
rect 123770 78618 124006 78854
rect 154490 78938 154726 79174
rect 154490 78618 154726 78854
rect 185210 78938 185446 79174
rect 185210 78618 185446 78854
rect 215930 78938 216166 79174
rect 215930 78618 216166 78854
rect 246650 78938 246886 79174
rect 246650 78618 246886 78854
rect 277370 78938 277606 79174
rect 277370 78618 277606 78854
rect 308090 78938 308326 79174
rect 308090 78618 308326 78854
rect 338810 78938 339046 79174
rect 338810 78618 339046 78854
rect 369530 78938 369766 79174
rect 369530 78618 369766 78854
rect 400250 78938 400486 79174
rect 400250 78618 400486 78854
rect 430970 78938 431206 79174
rect 430970 78618 431206 78854
rect 461690 78938 461926 79174
rect 461690 78618 461926 78854
rect 492410 78938 492646 79174
rect 492410 78618 492646 78854
rect 523130 78938 523366 79174
rect 523130 78618 523366 78854
rect 553850 78938 554086 79174
rect 553850 78618 554086 78854
rect 16250 75218 16486 75454
rect 16250 74898 16486 75134
rect 46970 75218 47206 75454
rect 46970 74898 47206 75134
rect 77690 75218 77926 75454
rect 77690 74898 77926 75134
rect 108410 75218 108646 75454
rect 108410 74898 108646 75134
rect 139130 75218 139366 75454
rect 139130 74898 139366 75134
rect 169850 75218 170086 75454
rect 169850 74898 170086 75134
rect 200570 75218 200806 75454
rect 200570 74898 200806 75134
rect 231290 75218 231526 75454
rect 231290 74898 231526 75134
rect 262010 75218 262246 75454
rect 262010 74898 262246 75134
rect 292730 75218 292966 75454
rect 292730 74898 292966 75134
rect 323450 75218 323686 75454
rect 323450 74898 323686 75134
rect 354170 75218 354406 75454
rect 354170 74898 354406 75134
rect 384890 75218 385126 75454
rect 384890 74898 385126 75134
rect 415610 75218 415846 75454
rect 415610 74898 415846 75134
rect 446330 75218 446566 75454
rect 446330 74898 446566 75134
rect 477050 75218 477286 75454
rect 477050 74898 477286 75134
rect 507770 75218 508006 75454
rect 507770 74898 508006 75134
rect 538490 75218 538726 75454
rect 538490 74898 538726 75134
rect 9266 46658 9502 46894
rect 9586 46658 9822 46894
rect 9266 46338 9502 46574
rect 9586 46338 9822 46574
rect 567866 65258 568102 65494
rect 568186 65258 568422 65494
rect 567866 64938 568102 65174
rect 568186 64938 568422 65174
rect 31610 42938 31846 43174
rect 31610 42618 31846 42854
rect 62330 42938 62566 43174
rect 62330 42618 62566 42854
rect 93050 42938 93286 43174
rect 93050 42618 93286 42854
rect 123770 42938 124006 43174
rect 123770 42618 124006 42854
rect 154490 42938 154726 43174
rect 154490 42618 154726 42854
rect 185210 42938 185446 43174
rect 185210 42618 185446 42854
rect 215930 42938 216166 43174
rect 215930 42618 216166 42854
rect 246650 42938 246886 43174
rect 246650 42618 246886 42854
rect 277370 42938 277606 43174
rect 277370 42618 277606 42854
rect 308090 42938 308326 43174
rect 308090 42618 308326 42854
rect 338810 42938 339046 43174
rect 338810 42618 339046 42854
rect 369530 42938 369766 43174
rect 369530 42618 369766 42854
rect 400250 42938 400486 43174
rect 400250 42618 400486 42854
rect 430970 42938 431206 43174
rect 430970 42618 431206 42854
rect 461690 42938 461926 43174
rect 461690 42618 461926 42854
rect 492410 42938 492646 43174
rect 492410 42618 492646 42854
rect 523130 42938 523366 43174
rect 523130 42618 523366 42854
rect 553850 42938 554086 43174
rect 553850 42618 554086 42854
rect 16250 39218 16486 39454
rect 16250 38898 16486 39134
rect 46970 39218 47206 39454
rect 46970 38898 47206 39134
rect 77690 39218 77926 39454
rect 77690 38898 77926 39134
rect 108410 39218 108646 39454
rect 108410 38898 108646 39134
rect 139130 39218 139366 39454
rect 139130 38898 139366 39134
rect 169850 39218 170086 39454
rect 169850 38898 170086 39134
rect 200570 39218 200806 39454
rect 200570 38898 200806 39134
rect 231290 39218 231526 39454
rect 231290 38898 231526 39134
rect 262010 39218 262246 39454
rect 262010 38898 262246 39134
rect 292730 39218 292966 39454
rect 292730 38898 292966 39134
rect 323450 39218 323686 39454
rect 323450 38898 323686 39134
rect 354170 39218 354406 39454
rect 354170 38898 354406 39134
rect 384890 39218 385126 39454
rect 384890 38898 385126 39134
rect 415610 39218 415846 39454
rect 415610 38898 415846 39134
rect 446330 39218 446566 39454
rect 446330 38898 446566 39134
rect 477050 39218 477286 39454
rect 477050 38898 477286 39134
rect 507770 39218 508006 39454
rect 507770 38898 508006 39134
rect 538490 39218 538726 39454
rect 538490 38898 538726 39134
rect 567866 29258 568102 29494
rect 568186 29258 568422 29494
rect 567866 28938 568102 29174
rect 568186 28938 568422 29174
rect 9266 10658 9502 10894
rect 9586 10658 9822 10894
rect 9266 10338 9502 10574
rect 9586 10338 9822 10574
rect 9266 -2502 9502 -2266
rect 9586 -2502 9822 -2266
rect 9266 -2822 9502 -2586
rect 9586 -2822 9822 -2586
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 41546 6938 41782 7174
rect 41866 6938 42102 7174
rect 41546 6618 41782 6854
rect 41866 6618 42102 6854
rect 41546 -1542 41782 -1306
rect 41866 -1542 42102 -1306
rect 41546 -1862 41782 -1626
rect 41866 -1862 42102 -1626
rect 45266 10658 45502 10894
rect 45586 10658 45822 10894
rect 45266 10338 45502 10574
rect 45586 10338 45822 10574
rect 45266 -2502 45502 -2266
rect 45586 -2502 45822 -2266
rect 45266 -2822 45502 -2586
rect 45586 -2822 45822 -2586
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 77546 6938 77782 7174
rect 77866 6938 78102 7174
rect 77546 6618 77782 6854
rect 77866 6618 78102 6854
rect 77546 -1542 77782 -1306
rect 77866 -1542 78102 -1306
rect 77546 -1862 77782 -1626
rect 77866 -1862 78102 -1626
rect 81266 10658 81502 10894
rect 81586 10658 81822 10894
rect 81266 10338 81502 10574
rect 81586 10338 81822 10574
rect 81266 -2502 81502 -2266
rect 81586 -2502 81822 -2266
rect 81266 -2822 81502 -2586
rect 81586 -2822 81822 -2586
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 113546 6938 113782 7174
rect 113866 6938 114102 7174
rect 113546 6618 113782 6854
rect 113866 6618 114102 6854
rect 113546 -1542 113782 -1306
rect 113866 -1542 114102 -1306
rect 113546 -1862 113782 -1626
rect 113866 -1862 114102 -1626
rect 117266 10658 117502 10894
rect 117586 10658 117822 10894
rect 117266 10338 117502 10574
rect 117586 10338 117822 10574
rect 117266 -2502 117502 -2266
rect 117586 -2502 117822 -2266
rect 117266 -2822 117502 -2586
rect 117586 -2822 117822 -2586
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 149546 6938 149782 7174
rect 149866 6938 150102 7174
rect 149546 6618 149782 6854
rect 149866 6618 150102 6854
rect 149546 -1542 149782 -1306
rect 149866 -1542 150102 -1306
rect 149546 -1862 149782 -1626
rect 149866 -1862 150102 -1626
rect 153266 10658 153502 10894
rect 153586 10658 153822 10894
rect 153266 10338 153502 10574
rect 153586 10338 153822 10574
rect 153266 -2502 153502 -2266
rect 153586 -2502 153822 -2266
rect 153266 -2822 153502 -2586
rect 153586 -2822 153822 -2586
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 185546 6938 185782 7174
rect 185866 6938 186102 7174
rect 185546 6618 185782 6854
rect 185866 6618 186102 6854
rect 185546 -1542 185782 -1306
rect 185866 -1542 186102 -1306
rect 185546 -1862 185782 -1626
rect 185866 -1862 186102 -1626
rect 189266 10658 189502 10894
rect 189586 10658 189822 10894
rect 189266 10338 189502 10574
rect 189586 10338 189822 10574
rect 189266 -2502 189502 -2266
rect 189586 -2502 189822 -2266
rect 189266 -2822 189502 -2586
rect 189586 -2822 189822 -2586
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 221546 6938 221782 7174
rect 221866 6938 222102 7174
rect 221546 6618 221782 6854
rect 221866 6618 222102 6854
rect 221546 -1542 221782 -1306
rect 221866 -1542 222102 -1306
rect 221546 -1862 221782 -1626
rect 221866 -1862 222102 -1626
rect 225266 10658 225502 10894
rect 225586 10658 225822 10894
rect 225266 10338 225502 10574
rect 225586 10338 225822 10574
rect 225266 -2502 225502 -2266
rect 225586 -2502 225822 -2266
rect 225266 -2822 225502 -2586
rect 225586 -2822 225822 -2586
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 257546 6938 257782 7174
rect 257866 6938 258102 7174
rect 257546 6618 257782 6854
rect 257866 6618 258102 6854
rect 257546 -1542 257782 -1306
rect 257866 -1542 258102 -1306
rect 257546 -1862 257782 -1626
rect 257866 -1862 258102 -1626
rect 261266 10658 261502 10894
rect 261586 10658 261822 10894
rect 261266 10338 261502 10574
rect 261586 10338 261822 10574
rect 261266 -2502 261502 -2266
rect 261586 -2502 261822 -2266
rect 261266 -2822 261502 -2586
rect 261586 -2822 261822 -2586
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 293546 6938 293782 7174
rect 293866 6938 294102 7174
rect 293546 6618 293782 6854
rect 293866 6618 294102 6854
rect 293546 -1542 293782 -1306
rect 293866 -1542 294102 -1306
rect 293546 -1862 293782 -1626
rect 293866 -1862 294102 -1626
rect 297266 10658 297502 10894
rect 297586 10658 297822 10894
rect 297266 10338 297502 10574
rect 297586 10338 297822 10574
rect 297266 -2502 297502 -2266
rect 297586 -2502 297822 -2266
rect 297266 -2822 297502 -2586
rect 297586 -2822 297822 -2586
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 329546 6938 329782 7174
rect 329866 6938 330102 7174
rect 329546 6618 329782 6854
rect 329866 6618 330102 6854
rect 329546 -1542 329782 -1306
rect 329866 -1542 330102 -1306
rect 329546 -1862 329782 -1626
rect 329866 -1862 330102 -1626
rect 333266 10658 333502 10894
rect 333586 10658 333822 10894
rect 333266 10338 333502 10574
rect 333586 10338 333822 10574
rect 333266 -2502 333502 -2266
rect 333586 -2502 333822 -2266
rect 333266 -2822 333502 -2586
rect 333586 -2822 333822 -2586
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 365546 6938 365782 7174
rect 365866 6938 366102 7174
rect 365546 6618 365782 6854
rect 365866 6618 366102 6854
rect 365546 -1542 365782 -1306
rect 365866 -1542 366102 -1306
rect 365546 -1862 365782 -1626
rect 365866 -1862 366102 -1626
rect 369266 10658 369502 10894
rect 369586 10658 369822 10894
rect 369266 10338 369502 10574
rect 369586 10338 369822 10574
rect 369266 -2502 369502 -2266
rect 369586 -2502 369822 -2266
rect 369266 -2822 369502 -2586
rect 369586 -2822 369822 -2586
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 401546 6938 401782 7174
rect 401866 6938 402102 7174
rect 401546 6618 401782 6854
rect 401866 6618 402102 6854
rect 401546 -1542 401782 -1306
rect 401866 -1542 402102 -1306
rect 401546 -1862 401782 -1626
rect 401866 -1862 402102 -1626
rect 405266 10658 405502 10894
rect 405586 10658 405822 10894
rect 405266 10338 405502 10574
rect 405586 10338 405822 10574
rect 405266 -2502 405502 -2266
rect 405586 -2502 405822 -2266
rect 405266 -2822 405502 -2586
rect 405586 -2822 405822 -2586
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 437546 6938 437782 7174
rect 437866 6938 438102 7174
rect 437546 6618 437782 6854
rect 437866 6618 438102 6854
rect 437546 -1542 437782 -1306
rect 437866 -1542 438102 -1306
rect 437546 -1862 437782 -1626
rect 437866 -1862 438102 -1626
rect 441266 10658 441502 10894
rect 441586 10658 441822 10894
rect 441266 10338 441502 10574
rect 441586 10338 441822 10574
rect 441266 -2502 441502 -2266
rect 441586 -2502 441822 -2266
rect 441266 -2822 441502 -2586
rect 441586 -2822 441822 -2586
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 473546 6938 473782 7174
rect 473866 6938 474102 7174
rect 473546 6618 473782 6854
rect 473866 6618 474102 6854
rect 473546 -1542 473782 -1306
rect 473866 -1542 474102 -1306
rect 473546 -1862 473782 -1626
rect 473866 -1862 474102 -1626
rect 477266 10658 477502 10894
rect 477586 10658 477822 10894
rect 477266 10338 477502 10574
rect 477586 10338 477822 10574
rect 477266 -2502 477502 -2266
rect 477586 -2502 477822 -2266
rect 477266 -2822 477502 -2586
rect 477586 -2822 477822 -2586
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 509546 6938 509782 7174
rect 509866 6938 510102 7174
rect 509546 6618 509782 6854
rect 509866 6618 510102 6854
rect 509546 -1542 509782 -1306
rect 509866 -1542 510102 -1306
rect 509546 -1862 509782 -1626
rect 509866 -1862 510102 -1626
rect 513266 10658 513502 10894
rect 513586 10658 513822 10894
rect 513266 10338 513502 10574
rect 513586 10338 513822 10574
rect 513266 -2502 513502 -2266
rect 513586 -2502 513822 -2266
rect 513266 -2822 513502 -2586
rect 513586 -2822 513822 -2586
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 545546 6938 545782 7174
rect 545866 6938 546102 7174
rect 545546 6618 545782 6854
rect 545866 6618 546102 6854
rect 545546 -1542 545782 -1306
rect 545866 -1542 546102 -1306
rect 545546 -1862 545782 -1626
rect 545866 -1862 546102 -1626
rect 549266 10658 549502 10894
rect 549586 10658 549822 10894
rect 549266 10338 549502 10574
rect 549586 10338 549822 10574
rect 549266 -2502 549502 -2266
rect 549586 -2502 549822 -2266
rect 549266 -2822 549502 -2586
rect 549586 -2822 549822 -2586
rect 567866 -7302 568102 -7066
rect 568186 -7302 568422 -7066
rect 567866 -7622 568102 -7386
rect 568186 -7622 568422 -7386
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 581546 705562 581782 705798
rect 581866 705562 582102 705798
rect 581546 705242 581782 705478
rect 581866 705242 582102 705478
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 581546 690938 581782 691174
rect 581866 690938 582102 691174
rect 581546 690618 581782 690854
rect 581866 690618 582102 690854
rect 581546 654938 581782 655174
rect 581866 654938 582102 655174
rect 581546 654618 581782 654854
rect 581866 654618 582102 654854
rect 581546 618938 581782 619174
rect 581866 618938 582102 619174
rect 581546 618618 581782 618854
rect 581866 618618 582102 618854
rect 581546 582938 581782 583174
rect 581866 582938 582102 583174
rect 581546 582618 581782 582854
rect 581866 582618 582102 582854
rect 581546 546938 581782 547174
rect 581866 546938 582102 547174
rect 581546 546618 581782 546854
rect 581866 546618 582102 546854
rect 581546 510938 581782 511174
rect 581866 510938 582102 511174
rect 581546 510618 581782 510854
rect 581866 510618 582102 510854
rect 581546 474938 581782 475174
rect 581866 474938 582102 475174
rect 581546 474618 581782 474854
rect 581866 474618 582102 474854
rect 581546 438938 581782 439174
rect 581866 438938 582102 439174
rect 581546 438618 581782 438854
rect 581866 438618 582102 438854
rect 581546 402938 581782 403174
rect 581866 402938 582102 403174
rect 581546 402618 581782 402854
rect 581866 402618 582102 402854
rect 581546 366938 581782 367174
rect 581866 366938 582102 367174
rect 581546 366618 581782 366854
rect 581866 366618 582102 366854
rect 581546 330938 581782 331174
rect 581866 330938 582102 331174
rect 581546 330618 581782 330854
rect 581866 330618 582102 330854
rect 581546 294938 581782 295174
rect 581866 294938 582102 295174
rect 581546 294618 581782 294854
rect 581866 294618 582102 294854
rect 581546 258938 581782 259174
rect 581866 258938 582102 259174
rect 581546 258618 581782 258854
rect 581866 258618 582102 258854
rect 581546 222938 581782 223174
rect 581866 222938 582102 223174
rect 581546 222618 581782 222854
rect 581866 222618 582102 222854
rect 581546 186938 581782 187174
rect 581866 186938 582102 187174
rect 581546 186618 581782 186854
rect 581866 186618 582102 186854
rect 581546 150938 581782 151174
rect 581866 150938 582102 151174
rect 581546 150618 581782 150854
rect 581866 150618 582102 150854
rect 581546 114938 581782 115174
rect 581866 114938 582102 115174
rect 581546 114618 581782 114854
rect 581866 114618 582102 114854
rect 581546 78938 581782 79174
rect 581866 78938 582102 79174
rect 581546 78618 581782 78854
rect 581866 78618 582102 78854
rect 581546 42938 581782 43174
rect 581866 42938 582102 43174
rect 581546 42618 581782 42854
rect 581866 42618 582102 42854
rect 581546 6938 581782 7174
rect 581866 6938 582102 7174
rect 581546 6618 581782 6854
rect 581866 6618 582102 6854
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 690938 586538 691174
rect 586622 690938 586858 691174
rect 586302 690618 586538 690854
rect 586622 690618 586858 690854
rect 586302 654938 586538 655174
rect 586622 654938 586858 655174
rect 586302 654618 586538 654854
rect 586622 654618 586858 654854
rect 586302 618938 586538 619174
rect 586622 618938 586858 619174
rect 586302 618618 586538 618854
rect 586622 618618 586858 618854
rect 586302 582938 586538 583174
rect 586622 582938 586858 583174
rect 586302 582618 586538 582854
rect 586622 582618 586858 582854
rect 586302 546938 586538 547174
rect 586622 546938 586858 547174
rect 586302 546618 586538 546854
rect 586622 546618 586858 546854
rect 586302 510938 586538 511174
rect 586622 510938 586858 511174
rect 586302 510618 586538 510854
rect 586622 510618 586858 510854
rect 586302 474938 586538 475174
rect 586622 474938 586858 475174
rect 586302 474618 586538 474854
rect 586622 474618 586858 474854
rect 586302 438938 586538 439174
rect 586622 438938 586858 439174
rect 586302 438618 586538 438854
rect 586622 438618 586858 438854
rect 586302 402938 586538 403174
rect 586622 402938 586858 403174
rect 586302 402618 586538 402854
rect 586622 402618 586858 402854
rect 586302 366938 586538 367174
rect 586622 366938 586858 367174
rect 586302 366618 586538 366854
rect 586622 366618 586858 366854
rect 586302 330938 586538 331174
rect 586622 330938 586858 331174
rect 586302 330618 586538 330854
rect 586622 330618 586858 330854
rect 586302 294938 586538 295174
rect 586622 294938 586858 295174
rect 586302 294618 586538 294854
rect 586622 294618 586858 294854
rect 586302 258938 586538 259174
rect 586622 258938 586858 259174
rect 586302 258618 586538 258854
rect 586622 258618 586858 258854
rect 586302 222938 586538 223174
rect 586622 222938 586858 223174
rect 586302 222618 586538 222854
rect 586622 222618 586858 222854
rect 586302 186938 586538 187174
rect 586622 186938 586858 187174
rect 586302 186618 586538 186854
rect 586622 186618 586858 186854
rect 586302 150938 586538 151174
rect 586622 150938 586858 151174
rect 586302 150618 586538 150854
rect 586622 150618 586858 150854
rect 586302 114938 586538 115174
rect 586622 114938 586858 115174
rect 586302 114618 586538 114854
rect 586622 114618 586858 114854
rect 586302 78938 586538 79174
rect 586622 78938 586858 79174
rect 586302 78618 586538 78854
rect 586622 78618 586858 78854
rect 586302 42938 586538 43174
rect 586622 42938 586858 43174
rect 586302 42618 586538 42854
rect 586622 42618 586858 42854
rect 586302 6938 586538 7174
rect 586622 6938 586858 7174
rect 586302 6618 586538 6854
rect 586622 6618 586858 6854
rect 581546 -1542 581782 -1306
rect 581866 -1542 582102 -1306
rect 581546 -1862 581782 -1626
rect 581866 -1862 582102 -1626
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 694658 587498 694894
rect 587582 694658 587818 694894
rect 587262 694338 587498 694574
rect 587582 694338 587818 694574
rect 587262 658658 587498 658894
rect 587582 658658 587818 658894
rect 587262 658338 587498 658574
rect 587582 658338 587818 658574
rect 587262 622658 587498 622894
rect 587582 622658 587818 622894
rect 587262 622338 587498 622574
rect 587582 622338 587818 622574
rect 587262 586658 587498 586894
rect 587582 586658 587818 586894
rect 587262 586338 587498 586574
rect 587582 586338 587818 586574
rect 587262 550658 587498 550894
rect 587582 550658 587818 550894
rect 587262 550338 587498 550574
rect 587582 550338 587818 550574
rect 587262 514658 587498 514894
rect 587582 514658 587818 514894
rect 587262 514338 587498 514574
rect 587582 514338 587818 514574
rect 587262 478658 587498 478894
rect 587582 478658 587818 478894
rect 587262 478338 587498 478574
rect 587582 478338 587818 478574
rect 587262 442658 587498 442894
rect 587582 442658 587818 442894
rect 587262 442338 587498 442574
rect 587582 442338 587818 442574
rect 587262 406658 587498 406894
rect 587582 406658 587818 406894
rect 587262 406338 587498 406574
rect 587582 406338 587818 406574
rect 587262 370658 587498 370894
rect 587582 370658 587818 370894
rect 587262 370338 587498 370574
rect 587582 370338 587818 370574
rect 587262 334658 587498 334894
rect 587582 334658 587818 334894
rect 587262 334338 587498 334574
rect 587582 334338 587818 334574
rect 587262 298658 587498 298894
rect 587582 298658 587818 298894
rect 587262 298338 587498 298574
rect 587582 298338 587818 298574
rect 587262 262658 587498 262894
rect 587582 262658 587818 262894
rect 587262 262338 587498 262574
rect 587582 262338 587818 262574
rect 587262 226658 587498 226894
rect 587582 226658 587818 226894
rect 587262 226338 587498 226574
rect 587582 226338 587818 226574
rect 587262 190658 587498 190894
rect 587582 190658 587818 190894
rect 587262 190338 587498 190574
rect 587582 190338 587818 190574
rect 587262 154658 587498 154894
rect 587582 154658 587818 154894
rect 587262 154338 587498 154574
rect 587582 154338 587818 154574
rect 587262 118658 587498 118894
rect 587582 118658 587818 118894
rect 587262 118338 587498 118574
rect 587582 118338 587818 118574
rect 587262 82658 587498 82894
rect 587582 82658 587818 82894
rect 587262 82338 587498 82574
rect 587582 82338 587818 82574
rect 587262 46658 587498 46894
rect 587582 46658 587818 46894
rect 587262 46338 587498 46574
rect 587582 46338 587818 46574
rect 587262 10658 587498 10894
rect 587582 10658 587818 10894
rect 587262 10338 587498 10574
rect 587582 10338 587818 10574
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 698378 588458 698614
rect 588542 698378 588778 698614
rect 588222 698058 588458 698294
rect 588542 698058 588778 698294
rect 588222 662378 588458 662614
rect 588542 662378 588778 662614
rect 588222 662058 588458 662294
rect 588542 662058 588778 662294
rect 588222 626378 588458 626614
rect 588542 626378 588778 626614
rect 588222 626058 588458 626294
rect 588542 626058 588778 626294
rect 588222 590378 588458 590614
rect 588542 590378 588778 590614
rect 588222 590058 588458 590294
rect 588542 590058 588778 590294
rect 588222 554378 588458 554614
rect 588542 554378 588778 554614
rect 588222 554058 588458 554294
rect 588542 554058 588778 554294
rect 588222 518378 588458 518614
rect 588542 518378 588778 518614
rect 588222 518058 588458 518294
rect 588542 518058 588778 518294
rect 588222 482378 588458 482614
rect 588542 482378 588778 482614
rect 588222 482058 588458 482294
rect 588542 482058 588778 482294
rect 588222 446378 588458 446614
rect 588542 446378 588778 446614
rect 588222 446058 588458 446294
rect 588542 446058 588778 446294
rect 588222 410378 588458 410614
rect 588542 410378 588778 410614
rect 588222 410058 588458 410294
rect 588542 410058 588778 410294
rect 588222 374378 588458 374614
rect 588542 374378 588778 374614
rect 588222 374058 588458 374294
rect 588542 374058 588778 374294
rect 588222 338378 588458 338614
rect 588542 338378 588778 338614
rect 588222 338058 588458 338294
rect 588542 338058 588778 338294
rect 588222 302378 588458 302614
rect 588542 302378 588778 302614
rect 588222 302058 588458 302294
rect 588542 302058 588778 302294
rect 588222 266378 588458 266614
rect 588542 266378 588778 266614
rect 588222 266058 588458 266294
rect 588542 266058 588778 266294
rect 588222 230378 588458 230614
rect 588542 230378 588778 230614
rect 588222 230058 588458 230294
rect 588542 230058 588778 230294
rect 588222 194378 588458 194614
rect 588542 194378 588778 194614
rect 588222 194058 588458 194294
rect 588542 194058 588778 194294
rect 588222 158378 588458 158614
rect 588542 158378 588778 158614
rect 588222 158058 588458 158294
rect 588542 158058 588778 158294
rect 588222 122378 588458 122614
rect 588542 122378 588778 122614
rect 588222 122058 588458 122294
rect 588542 122058 588778 122294
rect 588222 86378 588458 86614
rect 588542 86378 588778 86614
rect 588222 86058 588458 86294
rect 588542 86058 588778 86294
rect 588222 50378 588458 50614
rect 588542 50378 588778 50614
rect 588222 50058 588458 50294
rect 588542 50058 588778 50294
rect 588222 14378 588458 14614
rect 588542 14378 588778 14614
rect 588222 14058 588458 14294
rect 588542 14058 588778 14294
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 666098 589418 666334
rect 589502 666098 589738 666334
rect 589182 665778 589418 666014
rect 589502 665778 589738 666014
rect 589182 630098 589418 630334
rect 589502 630098 589738 630334
rect 589182 629778 589418 630014
rect 589502 629778 589738 630014
rect 589182 594098 589418 594334
rect 589502 594098 589738 594334
rect 589182 593778 589418 594014
rect 589502 593778 589738 594014
rect 589182 558098 589418 558334
rect 589502 558098 589738 558334
rect 589182 557778 589418 558014
rect 589502 557778 589738 558014
rect 589182 522098 589418 522334
rect 589502 522098 589738 522334
rect 589182 521778 589418 522014
rect 589502 521778 589738 522014
rect 589182 486098 589418 486334
rect 589502 486098 589738 486334
rect 589182 485778 589418 486014
rect 589502 485778 589738 486014
rect 589182 450098 589418 450334
rect 589502 450098 589738 450334
rect 589182 449778 589418 450014
rect 589502 449778 589738 450014
rect 589182 414098 589418 414334
rect 589502 414098 589738 414334
rect 589182 413778 589418 414014
rect 589502 413778 589738 414014
rect 589182 378098 589418 378334
rect 589502 378098 589738 378334
rect 589182 377778 589418 378014
rect 589502 377778 589738 378014
rect 589182 342098 589418 342334
rect 589502 342098 589738 342334
rect 589182 341778 589418 342014
rect 589502 341778 589738 342014
rect 589182 306098 589418 306334
rect 589502 306098 589738 306334
rect 589182 305778 589418 306014
rect 589502 305778 589738 306014
rect 589182 270098 589418 270334
rect 589502 270098 589738 270334
rect 589182 269778 589418 270014
rect 589502 269778 589738 270014
rect 589182 234098 589418 234334
rect 589502 234098 589738 234334
rect 589182 233778 589418 234014
rect 589502 233778 589738 234014
rect 589182 198098 589418 198334
rect 589502 198098 589738 198334
rect 589182 197778 589418 198014
rect 589502 197778 589738 198014
rect 589182 162098 589418 162334
rect 589502 162098 589738 162334
rect 589182 161778 589418 162014
rect 589502 161778 589738 162014
rect 589182 126098 589418 126334
rect 589502 126098 589738 126334
rect 589182 125778 589418 126014
rect 589502 125778 589738 126014
rect 589182 90098 589418 90334
rect 589502 90098 589738 90334
rect 589182 89778 589418 90014
rect 589502 89778 589738 90014
rect 589182 54098 589418 54334
rect 589502 54098 589738 54334
rect 589182 53778 589418 54014
rect 589502 53778 589738 54014
rect 589182 18098 589418 18334
rect 589502 18098 589738 18334
rect 589182 17778 589418 18014
rect 589502 17778 589738 18014
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 669818 590378 670054
rect 590462 669818 590698 670054
rect 590142 669498 590378 669734
rect 590462 669498 590698 669734
rect 590142 633818 590378 634054
rect 590462 633818 590698 634054
rect 590142 633498 590378 633734
rect 590462 633498 590698 633734
rect 590142 597818 590378 598054
rect 590462 597818 590698 598054
rect 590142 597498 590378 597734
rect 590462 597498 590698 597734
rect 590142 561818 590378 562054
rect 590462 561818 590698 562054
rect 590142 561498 590378 561734
rect 590462 561498 590698 561734
rect 590142 525818 590378 526054
rect 590462 525818 590698 526054
rect 590142 525498 590378 525734
rect 590462 525498 590698 525734
rect 590142 489818 590378 490054
rect 590462 489818 590698 490054
rect 590142 489498 590378 489734
rect 590462 489498 590698 489734
rect 590142 453818 590378 454054
rect 590462 453818 590698 454054
rect 590142 453498 590378 453734
rect 590462 453498 590698 453734
rect 590142 417818 590378 418054
rect 590462 417818 590698 418054
rect 590142 417498 590378 417734
rect 590462 417498 590698 417734
rect 590142 381818 590378 382054
rect 590462 381818 590698 382054
rect 590142 381498 590378 381734
rect 590462 381498 590698 381734
rect 590142 345818 590378 346054
rect 590462 345818 590698 346054
rect 590142 345498 590378 345734
rect 590462 345498 590698 345734
rect 590142 309818 590378 310054
rect 590462 309818 590698 310054
rect 590142 309498 590378 309734
rect 590462 309498 590698 309734
rect 590142 273818 590378 274054
rect 590462 273818 590698 274054
rect 590142 273498 590378 273734
rect 590462 273498 590698 273734
rect 590142 237818 590378 238054
rect 590462 237818 590698 238054
rect 590142 237498 590378 237734
rect 590462 237498 590698 237734
rect 590142 201818 590378 202054
rect 590462 201818 590698 202054
rect 590142 201498 590378 201734
rect 590462 201498 590698 201734
rect 590142 165818 590378 166054
rect 590462 165818 590698 166054
rect 590142 165498 590378 165734
rect 590462 165498 590698 165734
rect 590142 129818 590378 130054
rect 590462 129818 590698 130054
rect 590142 129498 590378 129734
rect 590462 129498 590698 129734
rect 590142 93818 590378 94054
rect 590462 93818 590698 94054
rect 590142 93498 590378 93734
rect 590462 93498 590698 93734
rect 590142 57818 590378 58054
rect 590462 57818 590698 58054
rect 590142 57498 590378 57734
rect 590462 57498 590698 57734
rect 590142 21818 590378 22054
rect 590462 21818 590698 22054
rect 590142 21498 590378 21734
rect 590462 21498 590698 21734
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 673538 591338 673774
rect 591422 673538 591658 673774
rect 591102 673218 591338 673454
rect 591422 673218 591658 673454
rect 591102 637538 591338 637774
rect 591422 637538 591658 637774
rect 591102 637218 591338 637454
rect 591422 637218 591658 637454
rect 591102 601538 591338 601774
rect 591422 601538 591658 601774
rect 591102 601218 591338 601454
rect 591422 601218 591658 601454
rect 591102 565538 591338 565774
rect 591422 565538 591658 565774
rect 591102 565218 591338 565454
rect 591422 565218 591658 565454
rect 591102 529538 591338 529774
rect 591422 529538 591658 529774
rect 591102 529218 591338 529454
rect 591422 529218 591658 529454
rect 591102 493538 591338 493774
rect 591422 493538 591658 493774
rect 591102 493218 591338 493454
rect 591422 493218 591658 493454
rect 591102 457538 591338 457774
rect 591422 457538 591658 457774
rect 591102 457218 591338 457454
rect 591422 457218 591658 457454
rect 591102 421538 591338 421774
rect 591422 421538 591658 421774
rect 591102 421218 591338 421454
rect 591422 421218 591658 421454
rect 591102 385538 591338 385774
rect 591422 385538 591658 385774
rect 591102 385218 591338 385454
rect 591422 385218 591658 385454
rect 591102 349538 591338 349774
rect 591422 349538 591658 349774
rect 591102 349218 591338 349454
rect 591422 349218 591658 349454
rect 591102 313538 591338 313774
rect 591422 313538 591658 313774
rect 591102 313218 591338 313454
rect 591422 313218 591658 313454
rect 591102 277538 591338 277774
rect 591422 277538 591658 277774
rect 591102 277218 591338 277454
rect 591422 277218 591658 277454
rect 591102 241538 591338 241774
rect 591422 241538 591658 241774
rect 591102 241218 591338 241454
rect 591422 241218 591658 241454
rect 591102 205538 591338 205774
rect 591422 205538 591658 205774
rect 591102 205218 591338 205454
rect 591422 205218 591658 205454
rect 591102 169538 591338 169774
rect 591422 169538 591658 169774
rect 591102 169218 591338 169454
rect 591422 169218 591658 169454
rect 591102 133538 591338 133774
rect 591422 133538 591658 133774
rect 591102 133218 591338 133454
rect 591422 133218 591658 133454
rect 591102 97538 591338 97774
rect 591422 97538 591658 97774
rect 591102 97218 591338 97454
rect 591422 97218 591658 97454
rect 591102 61538 591338 61774
rect 591422 61538 591658 61774
rect 591102 61218 591338 61454
rect 591422 61218 591658 61454
rect 591102 25538 591338 25774
rect 591422 25538 591658 25774
rect 591102 25218 591338 25454
rect 591422 25218 591658 25454
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 677258 592298 677494
rect 592382 677258 592618 677494
rect 592062 676938 592298 677174
rect 592382 676938 592618 677174
rect 592062 641258 592298 641494
rect 592382 641258 592618 641494
rect 592062 640938 592298 641174
rect 592382 640938 592618 641174
rect 592062 605258 592298 605494
rect 592382 605258 592618 605494
rect 592062 604938 592298 605174
rect 592382 604938 592618 605174
rect 592062 569258 592298 569494
rect 592382 569258 592618 569494
rect 592062 568938 592298 569174
rect 592382 568938 592618 569174
rect 592062 533258 592298 533494
rect 592382 533258 592618 533494
rect 592062 532938 592298 533174
rect 592382 532938 592618 533174
rect 592062 497258 592298 497494
rect 592382 497258 592618 497494
rect 592062 496938 592298 497174
rect 592382 496938 592618 497174
rect 592062 461258 592298 461494
rect 592382 461258 592618 461494
rect 592062 460938 592298 461174
rect 592382 460938 592618 461174
rect 592062 425258 592298 425494
rect 592382 425258 592618 425494
rect 592062 424938 592298 425174
rect 592382 424938 592618 425174
rect 592062 389258 592298 389494
rect 592382 389258 592618 389494
rect 592062 388938 592298 389174
rect 592382 388938 592618 389174
rect 592062 353258 592298 353494
rect 592382 353258 592618 353494
rect 592062 352938 592298 353174
rect 592382 352938 592618 353174
rect 592062 317258 592298 317494
rect 592382 317258 592618 317494
rect 592062 316938 592298 317174
rect 592382 316938 592618 317174
rect 592062 281258 592298 281494
rect 592382 281258 592618 281494
rect 592062 280938 592298 281174
rect 592382 280938 592618 281174
rect 592062 245258 592298 245494
rect 592382 245258 592618 245494
rect 592062 244938 592298 245174
rect 592382 244938 592618 245174
rect 592062 209258 592298 209494
rect 592382 209258 592618 209494
rect 592062 208938 592298 209174
rect 592382 208938 592618 209174
rect 592062 173258 592298 173494
rect 592382 173258 592618 173494
rect 592062 172938 592298 173174
rect 592382 172938 592618 173174
rect 592062 137258 592298 137494
rect 592382 137258 592618 137494
rect 592062 136938 592298 137174
rect 592382 136938 592618 137174
rect 592062 101258 592298 101494
rect 592382 101258 592618 101494
rect 592062 100938 592298 101174
rect 592382 100938 592618 101174
rect 592062 65258 592298 65494
rect 592382 65258 592618 65494
rect 592062 64938 592298 65174
rect 592382 64938 592618 65174
rect 592062 29258 592298 29494
rect 592382 29258 592618 29494
rect 592062 28938 592298 29174
rect 592382 28938 592618 29174
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 567866 711558
rect 568102 711322 568186 711558
rect 568422 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 567866 711238
rect 568102 711002 568186 711238
rect 568422 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 12986 707718
rect 13222 707482 13306 707718
rect 13542 707482 48986 707718
rect 49222 707482 49306 707718
rect 49542 707482 84986 707718
rect 85222 707482 85306 707718
rect 85542 707482 120986 707718
rect 121222 707482 121306 707718
rect 121542 707482 156986 707718
rect 157222 707482 157306 707718
rect 157542 707482 192986 707718
rect 193222 707482 193306 707718
rect 193542 707482 228986 707718
rect 229222 707482 229306 707718
rect 229542 707482 264986 707718
rect 265222 707482 265306 707718
rect 265542 707482 300986 707718
rect 301222 707482 301306 707718
rect 301542 707482 336986 707718
rect 337222 707482 337306 707718
rect 337542 707482 372986 707718
rect 373222 707482 373306 707718
rect 373542 707482 408986 707718
rect 409222 707482 409306 707718
rect 409542 707482 444986 707718
rect 445222 707482 445306 707718
rect 445542 707482 480986 707718
rect 481222 707482 481306 707718
rect 481542 707482 516986 707718
rect 517222 707482 517306 707718
rect 517542 707482 552986 707718
rect 553222 707482 553306 707718
rect 553542 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 12986 707398
rect 13222 707162 13306 707398
rect 13542 707162 48986 707398
rect 49222 707162 49306 707398
rect 49542 707162 84986 707398
rect 85222 707162 85306 707398
rect 85542 707162 120986 707398
rect 121222 707162 121306 707398
rect 121542 707162 156986 707398
rect 157222 707162 157306 707398
rect 157542 707162 192986 707398
rect 193222 707162 193306 707398
rect 193542 707162 228986 707398
rect 229222 707162 229306 707398
rect 229542 707162 264986 707398
rect 265222 707162 265306 707398
rect 265542 707162 300986 707398
rect 301222 707162 301306 707398
rect 301542 707162 336986 707398
rect 337222 707162 337306 707398
rect 337542 707162 372986 707398
rect 373222 707162 373306 707398
rect 373542 707162 408986 707398
rect 409222 707162 409306 707398
rect 409542 707162 444986 707398
rect 445222 707162 445306 707398
rect 445542 707162 480986 707398
rect 481222 707162 481306 707398
rect 481542 707162 516986 707398
rect 517222 707162 517306 707398
rect 517542 707162 552986 707398
rect 553222 707162 553306 707398
rect 553542 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 9266 706758
rect 9502 706522 9586 706758
rect 9822 706522 45266 706758
rect 45502 706522 45586 706758
rect 45822 706522 81266 706758
rect 81502 706522 81586 706758
rect 81822 706522 117266 706758
rect 117502 706522 117586 706758
rect 117822 706522 153266 706758
rect 153502 706522 153586 706758
rect 153822 706522 189266 706758
rect 189502 706522 189586 706758
rect 189822 706522 225266 706758
rect 225502 706522 225586 706758
rect 225822 706522 261266 706758
rect 261502 706522 261586 706758
rect 261822 706522 297266 706758
rect 297502 706522 297586 706758
rect 297822 706522 333266 706758
rect 333502 706522 333586 706758
rect 333822 706522 369266 706758
rect 369502 706522 369586 706758
rect 369822 706522 405266 706758
rect 405502 706522 405586 706758
rect 405822 706522 441266 706758
rect 441502 706522 441586 706758
rect 441822 706522 477266 706758
rect 477502 706522 477586 706758
rect 477822 706522 513266 706758
rect 513502 706522 513586 706758
rect 513822 706522 549266 706758
rect 549502 706522 549586 706758
rect 549822 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 9266 706438
rect 9502 706202 9586 706438
rect 9822 706202 45266 706438
rect 45502 706202 45586 706438
rect 45822 706202 81266 706438
rect 81502 706202 81586 706438
rect 81822 706202 117266 706438
rect 117502 706202 117586 706438
rect 117822 706202 153266 706438
rect 153502 706202 153586 706438
rect 153822 706202 189266 706438
rect 189502 706202 189586 706438
rect 189822 706202 225266 706438
rect 225502 706202 225586 706438
rect 225822 706202 261266 706438
rect 261502 706202 261586 706438
rect 261822 706202 297266 706438
rect 297502 706202 297586 706438
rect 297822 706202 333266 706438
rect 333502 706202 333586 706438
rect 333822 706202 369266 706438
rect 369502 706202 369586 706438
rect 369822 706202 405266 706438
rect 405502 706202 405586 706438
rect 405822 706202 441266 706438
rect 441502 706202 441586 706438
rect 441822 706202 477266 706438
rect 477502 706202 477586 706438
rect 477822 706202 513266 706438
rect 513502 706202 513586 706438
rect 513822 706202 549266 706438
rect 549502 706202 549586 706438
rect 549822 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 5546 705798
rect 5782 705562 5866 705798
rect 6102 705562 41546 705798
rect 41782 705562 41866 705798
rect 42102 705562 77546 705798
rect 77782 705562 77866 705798
rect 78102 705562 113546 705798
rect 113782 705562 113866 705798
rect 114102 705562 149546 705798
rect 149782 705562 149866 705798
rect 150102 705562 185546 705798
rect 185782 705562 185866 705798
rect 186102 705562 221546 705798
rect 221782 705562 221866 705798
rect 222102 705562 257546 705798
rect 257782 705562 257866 705798
rect 258102 705562 293546 705798
rect 293782 705562 293866 705798
rect 294102 705562 329546 705798
rect 329782 705562 329866 705798
rect 330102 705562 365546 705798
rect 365782 705562 365866 705798
rect 366102 705562 401546 705798
rect 401782 705562 401866 705798
rect 402102 705562 437546 705798
rect 437782 705562 437866 705798
rect 438102 705562 473546 705798
rect 473782 705562 473866 705798
rect 474102 705562 509546 705798
rect 509782 705562 509866 705798
rect 510102 705562 545546 705798
rect 545782 705562 545866 705798
rect 546102 705562 581546 705798
rect 581782 705562 581866 705798
rect 582102 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 5546 705478
rect 5782 705242 5866 705478
rect 6102 705242 41546 705478
rect 41782 705242 41866 705478
rect 42102 705242 77546 705478
rect 77782 705242 77866 705478
rect 78102 705242 113546 705478
rect 113782 705242 113866 705478
rect 114102 705242 149546 705478
rect 149782 705242 149866 705478
rect 150102 705242 185546 705478
rect 185782 705242 185866 705478
rect 186102 705242 221546 705478
rect 221782 705242 221866 705478
rect 222102 705242 257546 705478
rect 257782 705242 257866 705478
rect 258102 705242 293546 705478
rect 293782 705242 293866 705478
rect 294102 705242 329546 705478
rect 329782 705242 329866 705478
rect 330102 705242 365546 705478
rect 365782 705242 365866 705478
rect 366102 705242 401546 705478
rect 401782 705242 401866 705478
rect 402102 705242 437546 705478
rect 437782 705242 437866 705478
rect 438102 705242 473546 705478
rect 473782 705242 473866 705478
rect 474102 705242 509546 705478
rect 509782 705242 509866 705478
rect 510102 705242 545546 705478
rect 545782 705242 545866 705478
rect 546102 705242 581546 705478
rect 581782 705242 581866 705478
rect 582102 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 698614 592650 698646
rect -8726 698378 -4854 698614
rect -4618 698378 -4534 698614
rect -4298 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 588222 698614
rect 588458 698378 588542 698614
rect 588778 698378 592650 698614
rect -8726 698294 592650 698378
rect -8726 698058 -4854 698294
rect -4618 698058 -4534 698294
rect -4298 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 588222 698294
rect 588458 698058 588542 698294
rect 588778 698058 592650 698294
rect -8726 698026 592650 698058
rect -8726 694894 592650 694926
rect -8726 694658 -3894 694894
rect -3658 694658 -3574 694894
rect -3338 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 587262 694894
rect 587498 694658 587582 694894
rect 587818 694658 592650 694894
rect -8726 694574 592650 694658
rect -8726 694338 -3894 694574
rect -3658 694338 -3574 694574
rect -3338 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 587262 694574
rect 587498 694338 587582 694574
rect 587818 694338 592650 694574
rect -8726 694306 592650 694338
rect -8726 691174 592650 691206
rect -8726 690938 -2934 691174
rect -2698 690938 -2614 691174
rect -2378 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 586302 691174
rect 586538 690938 586622 691174
rect 586858 690938 592650 691174
rect -8726 690854 592650 690938
rect -8726 690618 -2934 690854
rect -2698 690618 -2614 690854
rect -2378 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 586302 690854
rect 586538 690618 586622 690854
rect 586858 690618 592650 690854
rect -8726 690586 592650 690618
rect -8726 687454 592650 687486
rect -8726 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 592650 687454
rect -8726 687134 592650 687218
rect -8726 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 592650 687134
rect -8726 686866 592650 686898
rect -8726 677494 592650 677526
rect -8726 677258 -8694 677494
rect -8458 677258 -8374 677494
rect -8138 677258 567866 677494
rect 568102 677258 568186 677494
rect 568422 677258 592062 677494
rect 592298 677258 592382 677494
rect 592618 677258 592650 677494
rect -8726 677174 592650 677258
rect -8726 676938 -8694 677174
rect -8458 676938 -8374 677174
rect -8138 676938 567866 677174
rect 568102 676938 568186 677174
rect 568422 676938 592062 677174
rect 592298 676938 592382 677174
rect 592618 676938 592650 677174
rect -8726 676906 592650 676938
rect -8726 673774 592650 673806
rect -8726 673538 -7734 673774
rect -7498 673538 -7414 673774
rect -7178 673538 591102 673774
rect 591338 673538 591422 673774
rect 591658 673538 592650 673774
rect -8726 673454 592650 673538
rect -8726 673218 -7734 673454
rect -7498 673218 -7414 673454
rect -7178 673218 591102 673454
rect 591338 673218 591422 673454
rect 591658 673218 592650 673454
rect -8726 673186 592650 673218
rect -8726 670054 592650 670086
rect -8726 669818 -6774 670054
rect -6538 669818 -6454 670054
rect -6218 669818 590142 670054
rect 590378 669818 590462 670054
rect 590698 669818 592650 670054
rect -8726 669734 592650 669818
rect -8726 669498 -6774 669734
rect -6538 669498 -6454 669734
rect -6218 669498 590142 669734
rect 590378 669498 590462 669734
rect 590698 669498 592650 669734
rect -8726 669466 592650 669498
rect -8726 666334 592650 666366
rect -8726 666098 -5814 666334
rect -5578 666098 -5494 666334
rect -5258 666098 589182 666334
rect 589418 666098 589502 666334
rect 589738 666098 592650 666334
rect -8726 666014 592650 666098
rect -8726 665778 -5814 666014
rect -5578 665778 -5494 666014
rect -5258 665778 589182 666014
rect 589418 665778 589502 666014
rect 589738 665778 592650 666014
rect -8726 665746 592650 665778
rect -8726 662614 592650 662646
rect -8726 662378 -4854 662614
rect -4618 662378 -4534 662614
rect -4298 662378 588222 662614
rect 588458 662378 588542 662614
rect 588778 662378 592650 662614
rect -8726 662294 592650 662378
rect -8726 662058 -4854 662294
rect -4618 662058 -4534 662294
rect -4298 662058 588222 662294
rect 588458 662058 588542 662294
rect 588778 662058 592650 662294
rect -8726 662026 592650 662058
rect -8726 658894 592650 658926
rect -8726 658658 -3894 658894
rect -3658 658658 -3574 658894
rect -3338 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 587262 658894
rect 587498 658658 587582 658894
rect 587818 658658 592650 658894
rect -8726 658574 592650 658658
rect -8726 658338 -3894 658574
rect -3658 658338 -3574 658574
rect -3338 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 587262 658574
rect 587498 658338 587582 658574
rect 587818 658338 592650 658574
rect -8726 658306 592650 658338
rect -8726 655174 592650 655206
rect -8726 654938 -2934 655174
rect -2698 654938 -2614 655174
rect -2378 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 31610 655174
rect 31846 654938 62330 655174
rect 62566 654938 93050 655174
rect 93286 654938 123770 655174
rect 124006 654938 154490 655174
rect 154726 654938 185210 655174
rect 185446 654938 215930 655174
rect 216166 654938 246650 655174
rect 246886 654938 277370 655174
rect 277606 654938 308090 655174
rect 308326 654938 338810 655174
rect 339046 654938 369530 655174
rect 369766 654938 400250 655174
rect 400486 654938 430970 655174
rect 431206 654938 461690 655174
rect 461926 654938 492410 655174
rect 492646 654938 523130 655174
rect 523366 654938 553850 655174
rect 554086 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 586302 655174
rect 586538 654938 586622 655174
rect 586858 654938 592650 655174
rect -8726 654854 592650 654938
rect -8726 654618 -2934 654854
rect -2698 654618 -2614 654854
rect -2378 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 31610 654854
rect 31846 654618 62330 654854
rect 62566 654618 93050 654854
rect 93286 654618 123770 654854
rect 124006 654618 154490 654854
rect 154726 654618 185210 654854
rect 185446 654618 215930 654854
rect 216166 654618 246650 654854
rect 246886 654618 277370 654854
rect 277606 654618 308090 654854
rect 308326 654618 338810 654854
rect 339046 654618 369530 654854
rect 369766 654618 400250 654854
rect 400486 654618 430970 654854
rect 431206 654618 461690 654854
rect 461926 654618 492410 654854
rect 492646 654618 523130 654854
rect 523366 654618 553850 654854
rect 554086 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 586302 654854
rect 586538 654618 586622 654854
rect 586858 654618 592650 654854
rect -8726 654586 592650 654618
rect -8726 651454 592650 651486
rect -8726 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 16250 651454
rect 16486 651218 46970 651454
rect 47206 651218 77690 651454
rect 77926 651218 108410 651454
rect 108646 651218 139130 651454
rect 139366 651218 169850 651454
rect 170086 651218 200570 651454
rect 200806 651218 231290 651454
rect 231526 651218 262010 651454
rect 262246 651218 292730 651454
rect 292966 651218 323450 651454
rect 323686 651218 354170 651454
rect 354406 651218 384890 651454
rect 385126 651218 415610 651454
rect 415846 651218 446330 651454
rect 446566 651218 477050 651454
rect 477286 651218 507770 651454
rect 508006 651218 538490 651454
rect 538726 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 592650 651454
rect -8726 651134 592650 651218
rect -8726 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 16250 651134
rect 16486 650898 46970 651134
rect 47206 650898 77690 651134
rect 77926 650898 108410 651134
rect 108646 650898 139130 651134
rect 139366 650898 169850 651134
rect 170086 650898 200570 651134
rect 200806 650898 231290 651134
rect 231526 650898 262010 651134
rect 262246 650898 292730 651134
rect 292966 650898 323450 651134
rect 323686 650898 354170 651134
rect 354406 650898 384890 651134
rect 385126 650898 415610 651134
rect 415846 650898 446330 651134
rect 446566 650898 477050 651134
rect 477286 650898 507770 651134
rect 508006 650898 538490 651134
rect 538726 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 592650 651134
rect -8726 650866 592650 650898
rect -8726 641494 592650 641526
rect -8726 641258 -8694 641494
rect -8458 641258 -8374 641494
rect -8138 641258 567866 641494
rect 568102 641258 568186 641494
rect 568422 641258 592062 641494
rect 592298 641258 592382 641494
rect 592618 641258 592650 641494
rect -8726 641174 592650 641258
rect -8726 640938 -8694 641174
rect -8458 640938 -8374 641174
rect -8138 640938 567866 641174
rect 568102 640938 568186 641174
rect 568422 640938 592062 641174
rect 592298 640938 592382 641174
rect 592618 640938 592650 641174
rect -8726 640906 592650 640938
rect -8726 637774 592650 637806
rect -8726 637538 -7734 637774
rect -7498 637538 -7414 637774
rect -7178 637538 591102 637774
rect 591338 637538 591422 637774
rect 591658 637538 592650 637774
rect -8726 637454 592650 637538
rect -8726 637218 -7734 637454
rect -7498 637218 -7414 637454
rect -7178 637218 591102 637454
rect 591338 637218 591422 637454
rect 591658 637218 592650 637454
rect -8726 637186 592650 637218
rect -8726 634054 592650 634086
rect -8726 633818 -6774 634054
rect -6538 633818 -6454 634054
rect -6218 633818 590142 634054
rect 590378 633818 590462 634054
rect 590698 633818 592650 634054
rect -8726 633734 592650 633818
rect -8726 633498 -6774 633734
rect -6538 633498 -6454 633734
rect -6218 633498 590142 633734
rect 590378 633498 590462 633734
rect 590698 633498 592650 633734
rect -8726 633466 592650 633498
rect -8726 630334 592650 630366
rect -8726 630098 -5814 630334
rect -5578 630098 -5494 630334
rect -5258 630098 589182 630334
rect 589418 630098 589502 630334
rect 589738 630098 592650 630334
rect -8726 630014 592650 630098
rect -8726 629778 -5814 630014
rect -5578 629778 -5494 630014
rect -5258 629778 589182 630014
rect 589418 629778 589502 630014
rect 589738 629778 592650 630014
rect -8726 629746 592650 629778
rect -8726 626614 592650 626646
rect -8726 626378 -4854 626614
rect -4618 626378 -4534 626614
rect -4298 626378 588222 626614
rect 588458 626378 588542 626614
rect 588778 626378 592650 626614
rect -8726 626294 592650 626378
rect -8726 626058 -4854 626294
rect -4618 626058 -4534 626294
rect -4298 626058 588222 626294
rect 588458 626058 588542 626294
rect 588778 626058 592650 626294
rect -8726 626026 592650 626058
rect -8726 622894 592650 622926
rect -8726 622658 -3894 622894
rect -3658 622658 -3574 622894
rect -3338 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 587262 622894
rect 587498 622658 587582 622894
rect 587818 622658 592650 622894
rect -8726 622574 592650 622658
rect -8726 622338 -3894 622574
rect -3658 622338 -3574 622574
rect -3338 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 587262 622574
rect 587498 622338 587582 622574
rect 587818 622338 592650 622574
rect -8726 622306 592650 622338
rect -8726 619174 592650 619206
rect -8726 618938 -2934 619174
rect -2698 618938 -2614 619174
rect -2378 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 31610 619174
rect 31846 618938 62330 619174
rect 62566 618938 93050 619174
rect 93286 618938 123770 619174
rect 124006 618938 154490 619174
rect 154726 618938 185210 619174
rect 185446 618938 215930 619174
rect 216166 618938 246650 619174
rect 246886 618938 277370 619174
rect 277606 618938 308090 619174
rect 308326 618938 338810 619174
rect 339046 618938 369530 619174
rect 369766 618938 400250 619174
rect 400486 618938 430970 619174
rect 431206 618938 461690 619174
rect 461926 618938 492410 619174
rect 492646 618938 523130 619174
rect 523366 618938 553850 619174
rect 554086 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 586302 619174
rect 586538 618938 586622 619174
rect 586858 618938 592650 619174
rect -8726 618854 592650 618938
rect -8726 618618 -2934 618854
rect -2698 618618 -2614 618854
rect -2378 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 31610 618854
rect 31846 618618 62330 618854
rect 62566 618618 93050 618854
rect 93286 618618 123770 618854
rect 124006 618618 154490 618854
rect 154726 618618 185210 618854
rect 185446 618618 215930 618854
rect 216166 618618 246650 618854
rect 246886 618618 277370 618854
rect 277606 618618 308090 618854
rect 308326 618618 338810 618854
rect 339046 618618 369530 618854
rect 369766 618618 400250 618854
rect 400486 618618 430970 618854
rect 431206 618618 461690 618854
rect 461926 618618 492410 618854
rect 492646 618618 523130 618854
rect 523366 618618 553850 618854
rect 554086 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 586302 618854
rect 586538 618618 586622 618854
rect 586858 618618 592650 618854
rect -8726 618586 592650 618618
rect -8726 615454 592650 615486
rect -8726 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 16250 615454
rect 16486 615218 46970 615454
rect 47206 615218 77690 615454
rect 77926 615218 108410 615454
rect 108646 615218 139130 615454
rect 139366 615218 169850 615454
rect 170086 615218 200570 615454
rect 200806 615218 231290 615454
rect 231526 615218 262010 615454
rect 262246 615218 292730 615454
rect 292966 615218 323450 615454
rect 323686 615218 354170 615454
rect 354406 615218 384890 615454
rect 385126 615218 415610 615454
rect 415846 615218 446330 615454
rect 446566 615218 477050 615454
rect 477286 615218 507770 615454
rect 508006 615218 538490 615454
rect 538726 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 592650 615454
rect -8726 615134 592650 615218
rect -8726 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 16250 615134
rect 16486 614898 46970 615134
rect 47206 614898 77690 615134
rect 77926 614898 108410 615134
rect 108646 614898 139130 615134
rect 139366 614898 169850 615134
rect 170086 614898 200570 615134
rect 200806 614898 231290 615134
rect 231526 614898 262010 615134
rect 262246 614898 292730 615134
rect 292966 614898 323450 615134
rect 323686 614898 354170 615134
rect 354406 614898 384890 615134
rect 385126 614898 415610 615134
rect 415846 614898 446330 615134
rect 446566 614898 477050 615134
rect 477286 614898 507770 615134
rect 508006 614898 538490 615134
rect 538726 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 592650 615134
rect -8726 614866 592650 614898
rect -8726 605494 592650 605526
rect -8726 605258 -8694 605494
rect -8458 605258 -8374 605494
rect -8138 605258 567866 605494
rect 568102 605258 568186 605494
rect 568422 605258 592062 605494
rect 592298 605258 592382 605494
rect 592618 605258 592650 605494
rect -8726 605174 592650 605258
rect -8726 604938 -8694 605174
rect -8458 604938 -8374 605174
rect -8138 604938 567866 605174
rect 568102 604938 568186 605174
rect 568422 604938 592062 605174
rect 592298 604938 592382 605174
rect 592618 604938 592650 605174
rect -8726 604906 592650 604938
rect -8726 601774 592650 601806
rect -8726 601538 -7734 601774
rect -7498 601538 -7414 601774
rect -7178 601538 591102 601774
rect 591338 601538 591422 601774
rect 591658 601538 592650 601774
rect -8726 601454 592650 601538
rect -8726 601218 -7734 601454
rect -7498 601218 -7414 601454
rect -7178 601218 591102 601454
rect 591338 601218 591422 601454
rect 591658 601218 592650 601454
rect -8726 601186 592650 601218
rect -8726 598054 592650 598086
rect -8726 597818 -6774 598054
rect -6538 597818 -6454 598054
rect -6218 597818 590142 598054
rect 590378 597818 590462 598054
rect 590698 597818 592650 598054
rect -8726 597734 592650 597818
rect -8726 597498 -6774 597734
rect -6538 597498 -6454 597734
rect -6218 597498 590142 597734
rect 590378 597498 590462 597734
rect 590698 597498 592650 597734
rect -8726 597466 592650 597498
rect -8726 594334 592650 594366
rect -8726 594098 -5814 594334
rect -5578 594098 -5494 594334
rect -5258 594098 589182 594334
rect 589418 594098 589502 594334
rect 589738 594098 592650 594334
rect -8726 594014 592650 594098
rect -8726 593778 -5814 594014
rect -5578 593778 -5494 594014
rect -5258 593778 589182 594014
rect 589418 593778 589502 594014
rect 589738 593778 592650 594014
rect -8726 593746 592650 593778
rect -8726 590614 592650 590646
rect -8726 590378 -4854 590614
rect -4618 590378 -4534 590614
rect -4298 590378 588222 590614
rect 588458 590378 588542 590614
rect 588778 590378 592650 590614
rect -8726 590294 592650 590378
rect -8726 590058 -4854 590294
rect -4618 590058 -4534 590294
rect -4298 590058 588222 590294
rect 588458 590058 588542 590294
rect 588778 590058 592650 590294
rect -8726 590026 592650 590058
rect -8726 586894 592650 586926
rect -8726 586658 -3894 586894
rect -3658 586658 -3574 586894
rect -3338 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 587262 586894
rect 587498 586658 587582 586894
rect 587818 586658 592650 586894
rect -8726 586574 592650 586658
rect -8726 586338 -3894 586574
rect -3658 586338 -3574 586574
rect -3338 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 587262 586574
rect 587498 586338 587582 586574
rect 587818 586338 592650 586574
rect -8726 586306 592650 586338
rect -8726 583174 592650 583206
rect -8726 582938 -2934 583174
rect -2698 582938 -2614 583174
rect -2378 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 31610 583174
rect 31846 582938 62330 583174
rect 62566 582938 93050 583174
rect 93286 582938 123770 583174
rect 124006 582938 154490 583174
rect 154726 582938 185210 583174
rect 185446 582938 215930 583174
rect 216166 582938 246650 583174
rect 246886 582938 277370 583174
rect 277606 582938 308090 583174
rect 308326 582938 338810 583174
rect 339046 582938 369530 583174
rect 369766 582938 400250 583174
rect 400486 582938 430970 583174
rect 431206 582938 461690 583174
rect 461926 582938 492410 583174
rect 492646 582938 523130 583174
rect 523366 582938 553850 583174
rect 554086 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 586302 583174
rect 586538 582938 586622 583174
rect 586858 582938 592650 583174
rect -8726 582854 592650 582938
rect -8726 582618 -2934 582854
rect -2698 582618 -2614 582854
rect -2378 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 31610 582854
rect 31846 582618 62330 582854
rect 62566 582618 93050 582854
rect 93286 582618 123770 582854
rect 124006 582618 154490 582854
rect 154726 582618 185210 582854
rect 185446 582618 215930 582854
rect 216166 582618 246650 582854
rect 246886 582618 277370 582854
rect 277606 582618 308090 582854
rect 308326 582618 338810 582854
rect 339046 582618 369530 582854
rect 369766 582618 400250 582854
rect 400486 582618 430970 582854
rect 431206 582618 461690 582854
rect 461926 582618 492410 582854
rect 492646 582618 523130 582854
rect 523366 582618 553850 582854
rect 554086 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 586302 582854
rect 586538 582618 586622 582854
rect 586858 582618 592650 582854
rect -8726 582586 592650 582618
rect -8726 579454 592650 579486
rect -8726 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 16250 579454
rect 16486 579218 46970 579454
rect 47206 579218 77690 579454
rect 77926 579218 108410 579454
rect 108646 579218 139130 579454
rect 139366 579218 169850 579454
rect 170086 579218 200570 579454
rect 200806 579218 231290 579454
rect 231526 579218 262010 579454
rect 262246 579218 292730 579454
rect 292966 579218 323450 579454
rect 323686 579218 354170 579454
rect 354406 579218 384890 579454
rect 385126 579218 415610 579454
rect 415846 579218 446330 579454
rect 446566 579218 477050 579454
rect 477286 579218 507770 579454
rect 508006 579218 538490 579454
rect 538726 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 592650 579454
rect -8726 579134 592650 579218
rect -8726 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 16250 579134
rect 16486 578898 46970 579134
rect 47206 578898 77690 579134
rect 77926 578898 108410 579134
rect 108646 578898 139130 579134
rect 139366 578898 169850 579134
rect 170086 578898 200570 579134
rect 200806 578898 231290 579134
rect 231526 578898 262010 579134
rect 262246 578898 292730 579134
rect 292966 578898 323450 579134
rect 323686 578898 354170 579134
rect 354406 578898 384890 579134
rect 385126 578898 415610 579134
rect 415846 578898 446330 579134
rect 446566 578898 477050 579134
rect 477286 578898 507770 579134
rect 508006 578898 538490 579134
rect 538726 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 592650 579134
rect -8726 578866 592650 578898
rect -8726 569494 592650 569526
rect -8726 569258 -8694 569494
rect -8458 569258 -8374 569494
rect -8138 569258 567866 569494
rect 568102 569258 568186 569494
rect 568422 569258 592062 569494
rect 592298 569258 592382 569494
rect 592618 569258 592650 569494
rect -8726 569174 592650 569258
rect -8726 568938 -8694 569174
rect -8458 568938 -8374 569174
rect -8138 568938 567866 569174
rect 568102 568938 568186 569174
rect 568422 568938 592062 569174
rect 592298 568938 592382 569174
rect 592618 568938 592650 569174
rect -8726 568906 592650 568938
rect -8726 565774 592650 565806
rect -8726 565538 -7734 565774
rect -7498 565538 -7414 565774
rect -7178 565538 591102 565774
rect 591338 565538 591422 565774
rect 591658 565538 592650 565774
rect -8726 565454 592650 565538
rect -8726 565218 -7734 565454
rect -7498 565218 -7414 565454
rect -7178 565218 591102 565454
rect 591338 565218 591422 565454
rect 591658 565218 592650 565454
rect -8726 565186 592650 565218
rect -8726 562054 592650 562086
rect -8726 561818 -6774 562054
rect -6538 561818 -6454 562054
rect -6218 561818 590142 562054
rect 590378 561818 590462 562054
rect 590698 561818 592650 562054
rect -8726 561734 592650 561818
rect -8726 561498 -6774 561734
rect -6538 561498 -6454 561734
rect -6218 561498 590142 561734
rect 590378 561498 590462 561734
rect 590698 561498 592650 561734
rect -8726 561466 592650 561498
rect -8726 558334 592650 558366
rect -8726 558098 -5814 558334
rect -5578 558098 -5494 558334
rect -5258 558098 589182 558334
rect 589418 558098 589502 558334
rect 589738 558098 592650 558334
rect -8726 558014 592650 558098
rect -8726 557778 -5814 558014
rect -5578 557778 -5494 558014
rect -5258 557778 589182 558014
rect 589418 557778 589502 558014
rect 589738 557778 592650 558014
rect -8726 557746 592650 557778
rect -8726 554614 592650 554646
rect -8726 554378 -4854 554614
rect -4618 554378 -4534 554614
rect -4298 554378 588222 554614
rect 588458 554378 588542 554614
rect 588778 554378 592650 554614
rect -8726 554294 592650 554378
rect -8726 554058 -4854 554294
rect -4618 554058 -4534 554294
rect -4298 554058 588222 554294
rect 588458 554058 588542 554294
rect 588778 554058 592650 554294
rect -8726 554026 592650 554058
rect -8726 550894 592650 550926
rect -8726 550658 -3894 550894
rect -3658 550658 -3574 550894
rect -3338 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 587262 550894
rect 587498 550658 587582 550894
rect 587818 550658 592650 550894
rect -8726 550574 592650 550658
rect -8726 550338 -3894 550574
rect -3658 550338 -3574 550574
rect -3338 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 587262 550574
rect 587498 550338 587582 550574
rect 587818 550338 592650 550574
rect -8726 550306 592650 550338
rect -8726 547174 592650 547206
rect -8726 546938 -2934 547174
rect -2698 546938 -2614 547174
rect -2378 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 31610 547174
rect 31846 546938 62330 547174
rect 62566 546938 93050 547174
rect 93286 546938 123770 547174
rect 124006 546938 154490 547174
rect 154726 546938 185210 547174
rect 185446 546938 215930 547174
rect 216166 546938 246650 547174
rect 246886 546938 277370 547174
rect 277606 546938 308090 547174
rect 308326 546938 338810 547174
rect 339046 546938 369530 547174
rect 369766 546938 400250 547174
rect 400486 546938 430970 547174
rect 431206 546938 461690 547174
rect 461926 546938 492410 547174
rect 492646 546938 523130 547174
rect 523366 546938 553850 547174
rect 554086 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 586302 547174
rect 586538 546938 586622 547174
rect 586858 546938 592650 547174
rect -8726 546854 592650 546938
rect -8726 546618 -2934 546854
rect -2698 546618 -2614 546854
rect -2378 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 31610 546854
rect 31846 546618 62330 546854
rect 62566 546618 93050 546854
rect 93286 546618 123770 546854
rect 124006 546618 154490 546854
rect 154726 546618 185210 546854
rect 185446 546618 215930 546854
rect 216166 546618 246650 546854
rect 246886 546618 277370 546854
rect 277606 546618 308090 546854
rect 308326 546618 338810 546854
rect 339046 546618 369530 546854
rect 369766 546618 400250 546854
rect 400486 546618 430970 546854
rect 431206 546618 461690 546854
rect 461926 546618 492410 546854
rect 492646 546618 523130 546854
rect 523366 546618 553850 546854
rect 554086 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 586302 546854
rect 586538 546618 586622 546854
rect 586858 546618 592650 546854
rect -8726 546586 592650 546618
rect -8726 543454 592650 543486
rect -8726 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 16250 543454
rect 16486 543218 46970 543454
rect 47206 543218 77690 543454
rect 77926 543218 108410 543454
rect 108646 543218 139130 543454
rect 139366 543218 169850 543454
rect 170086 543218 200570 543454
rect 200806 543218 231290 543454
rect 231526 543218 262010 543454
rect 262246 543218 292730 543454
rect 292966 543218 323450 543454
rect 323686 543218 354170 543454
rect 354406 543218 384890 543454
rect 385126 543218 415610 543454
rect 415846 543218 446330 543454
rect 446566 543218 477050 543454
rect 477286 543218 507770 543454
rect 508006 543218 538490 543454
rect 538726 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 592650 543454
rect -8726 543134 592650 543218
rect -8726 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 16250 543134
rect 16486 542898 46970 543134
rect 47206 542898 77690 543134
rect 77926 542898 108410 543134
rect 108646 542898 139130 543134
rect 139366 542898 169850 543134
rect 170086 542898 200570 543134
rect 200806 542898 231290 543134
rect 231526 542898 262010 543134
rect 262246 542898 292730 543134
rect 292966 542898 323450 543134
rect 323686 542898 354170 543134
rect 354406 542898 384890 543134
rect 385126 542898 415610 543134
rect 415846 542898 446330 543134
rect 446566 542898 477050 543134
rect 477286 542898 507770 543134
rect 508006 542898 538490 543134
rect 538726 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 592650 543134
rect -8726 542866 592650 542898
rect -8726 533494 592650 533526
rect -8726 533258 -8694 533494
rect -8458 533258 -8374 533494
rect -8138 533258 567866 533494
rect 568102 533258 568186 533494
rect 568422 533258 592062 533494
rect 592298 533258 592382 533494
rect 592618 533258 592650 533494
rect -8726 533174 592650 533258
rect -8726 532938 -8694 533174
rect -8458 532938 -8374 533174
rect -8138 532938 567866 533174
rect 568102 532938 568186 533174
rect 568422 532938 592062 533174
rect 592298 532938 592382 533174
rect 592618 532938 592650 533174
rect -8726 532906 592650 532938
rect -8726 529774 592650 529806
rect -8726 529538 -7734 529774
rect -7498 529538 -7414 529774
rect -7178 529538 591102 529774
rect 591338 529538 591422 529774
rect 591658 529538 592650 529774
rect -8726 529454 592650 529538
rect -8726 529218 -7734 529454
rect -7498 529218 -7414 529454
rect -7178 529218 591102 529454
rect 591338 529218 591422 529454
rect 591658 529218 592650 529454
rect -8726 529186 592650 529218
rect -8726 526054 592650 526086
rect -8726 525818 -6774 526054
rect -6538 525818 -6454 526054
rect -6218 525818 590142 526054
rect 590378 525818 590462 526054
rect 590698 525818 592650 526054
rect -8726 525734 592650 525818
rect -8726 525498 -6774 525734
rect -6538 525498 -6454 525734
rect -6218 525498 590142 525734
rect 590378 525498 590462 525734
rect 590698 525498 592650 525734
rect -8726 525466 592650 525498
rect -8726 522334 592650 522366
rect -8726 522098 -5814 522334
rect -5578 522098 -5494 522334
rect -5258 522098 589182 522334
rect 589418 522098 589502 522334
rect 589738 522098 592650 522334
rect -8726 522014 592650 522098
rect -8726 521778 -5814 522014
rect -5578 521778 -5494 522014
rect -5258 521778 589182 522014
rect 589418 521778 589502 522014
rect 589738 521778 592650 522014
rect -8726 521746 592650 521778
rect -8726 518614 592650 518646
rect -8726 518378 -4854 518614
rect -4618 518378 -4534 518614
rect -4298 518378 588222 518614
rect 588458 518378 588542 518614
rect 588778 518378 592650 518614
rect -8726 518294 592650 518378
rect -8726 518058 -4854 518294
rect -4618 518058 -4534 518294
rect -4298 518058 588222 518294
rect 588458 518058 588542 518294
rect 588778 518058 592650 518294
rect -8726 518026 592650 518058
rect -8726 514894 592650 514926
rect -8726 514658 -3894 514894
rect -3658 514658 -3574 514894
rect -3338 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 587262 514894
rect 587498 514658 587582 514894
rect 587818 514658 592650 514894
rect -8726 514574 592650 514658
rect -8726 514338 -3894 514574
rect -3658 514338 -3574 514574
rect -3338 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 587262 514574
rect 587498 514338 587582 514574
rect 587818 514338 592650 514574
rect -8726 514306 592650 514338
rect -8726 511174 592650 511206
rect -8726 510938 -2934 511174
rect -2698 510938 -2614 511174
rect -2378 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 31610 511174
rect 31846 510938 62330 511174
rect 62566 510938 93050 511174
rect 93286 510938 123770 511174
rect 124006 510938 154490 511174
rect 154726 510938 185210 511174
rect 185446 510938 215930 511174
rect 216166 510938 246650 511174
rect 246886 510938 277370 511174
rect 277606 510938 308090 511174
rect 308326 510938 338810 511174
rect 339046 510938 369530 511174
rect 369766 510938 400250 511174
rect 400486 510938 430970 511174
rect 431206 510938 461690 511174
rect 461926 510938 492410 511174
rect 492646 510938 523130 511174
rect 523366 510938 553850 511174
rect 554086 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 586302 511174
rect 586538 510938 586622 511174
rect 586858 510938 592650 511174
rect -8726 510854 592650 510938
rect -8726 510618 -2934 510854
rect -2698 510618 -2614 510854
rect -2378 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 31610 510854
rect 31846 510618 62330 510854
rect 62566 510618 93050 510854
rect 93286 510618 123770 510854
rect 124006 510618 154490 510854
rect 154726 510618 185210 510854
rect 185446 510618 215930 510854
rect 216166 510618 246650 510854
rect 246886 510618 277370 510854
rect 277606 510618 308090 510854
rect 308326 510618 338810 510854
rect 339046 510618 369530 510854
rect 369766 510618 400250 510854
rect 400486 510618 430970 510854
rect 431206 510618 461690 510854
rect 461926 510618 492410 510854
rect 492646 510618 523130 510854
rect 523366 510618 553850 510854
rect 554086 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 586302 510854
rect 586538 510618 586622 510854
rect 586858 510618 592650 510854
rect -8726 510586 592650 510618
rect -8726 507454 592650 507486
rect -8726 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 16250 507454
rect 16486 507218 46970 507454
rect 47206 507218 77690 507454
rect 77926 507218 108410 507454
rect 108646 507218 139130 507454
rect 139366 507218 169850 507454
rect 170086 507218 200570 507454
rect 200806 507218 231290 507454
rect 231526 507218 262010 507454
rect 262246 507218 292730 507454
rect 292966 507218 323450 507454
rect 323686 507218 354170 507454
rect 354406 507218 384890 507454
rect 385126 507218 415610 507454
rect 415846 507218 446330 507454
rect 446566 507218 477050 507454
rect 477286 507218 507770 507454
rect 508006 507218 538490 507454
rect 538726 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 592650 507454
rect -8726 507134 592650 507218
rect -8726 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 16250 507134
rect 16486 506898 46970 507134
rect 47206 506898 77690 507134
rect 77926 506898 108410 507134
rect 108646 506898 139130 507134
rect 139366 506898 169850 507134
rect 170086 506898 200570 507134
rect 200806 506898 231290 507134
rect 231526 506898 262010 507134
rect 262246 506898 292730 507134
rect 292966 506898 323450 507134
rect 323686 506898 354170 507134
rect 354406 506898 384890 507134
rect 385126 506898 415610 507134
rect 415846 506898 446330 507134
rect 446566 506898 477050 507134
rect 477286 506898 507770 507134
rect 508006 506898 538490 507134
rect 538726 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 592650 507134
rect -8726 506866 592650 506898
rect -8726 497494 592650 497526
rect -8726 497258 -8694 497494
rect -8458 497258 -8374 497494
rect -8138 497258 567866 497494
rect 568102 497258 568186 497494
rect 568422 497258 592062 497494
rect 592298 497258 592382 497494
rect 592618 497258 592650 497494
rect -8726 497174 592650 497258
rect -8726 496938 -8694 497174
rect -8458 496938 -8374 497174
rect -8138 496938 567866 497174
rect 568102 496938 568186 497174
rect 568422 496938 592062 497174
rect 592298 496938 592382 497174
rect 592618 496938 592650 497174
rect -8726 496906 592650 496938
rect -8726 493774 592650 493806
rect -8726 493538 -7734 493774
rect -7498 493538 -7414 493774
rect -7178 493538 591102 493774
rect 591338 493538 591422 493774
rect 591658 493538 592650 493774
rect -8726 493454 592650 493538
rect -8726 493218 -7734 493454
rect -7498 493218 -7414 493454
rect -7178 493218 591102 493454
rect 591338 493218 591422 493454
rect 591658 493218 592650 493454
rect -8726 493186 592650 493218
rect -8726 490054 592650 490086
rect -8726 489818 -6774 490054
rect -6538 489818 -6454 490054
rect -6218 489818 590142 490054
rect 590378 489818 590462 490054
rect 590698 489818 592650 490054
rect -8726 489734 592650 489818
rect -8726 489498 -6774 489734
rect -6538 489498 -6454 489734
rect -6218 489498 590142 489734
rect 590378 489498 590462 489734
rect 590698 489498 592650 489734
rect -8726 489466 592650 489498
rect -8726 486334 592650 486366
rect -8726 486098 -5814 486334
rect -5578 486098 -5494 486334
rect -5258 486098 589182 486334
rect 589418 486098 589502 486334
rect 589738 486098 592650 486334
rect -8726 486014 592650 486098
rect -8726 485778 -5814 486014
rect -5578 485778 -5494 486014
rect -5258 485778 589182 486014
rect 589418 485778 589502 486014
rect 589738 485778 592650 486014
rect -8726 485746 592650 485778
rect -8726 482614 592650 482646
rect -8726 482378 -4854 482614
rect -4618 482378 -4534 482614
rect -4298 482378 588222 482614
rect 588458 482378 588542 482614
rect 588778 482378 592650 482614
rect -8726 482294 592650 482378
rect -8726 482058 -4854 482294
rect -4618 482058 -4534 482294
rect -4298 482058 588222 482294
rect 588458 482058 588542 482294
rect 588778 482058 592650 482294
rect -8726 482026 592650 482058
rect -8726 478894 592650 478926
rect -8726 478658 -3894 478894
rect -3658 478658 -3574 478894
rect -3338 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 587262 478894
rect 587498 478658 587582 478894
rect 587818 478658 592650 478894
rect -8726 478574 592650 478658
rect -8726 478338 -3894 478574
rect -3658 478338 -3574 478574
rect -3338 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 587262 478574
rect 587498 478338 587582 478574
rect 587818 478338 592650 478574
rect -8726 478306 592650 478338
rect -8726 475174 592650 475206
rect -8726 474938 -2934 475174
rect -2698 474938 -2614 475174
rect -2378 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 31610 475174
rect 31846 474938 62330 475174
rect 62566 474938 93050 475174
rect 93286 474938 123770 475174
rect 124006 474938 154490 475174
rect 154726 474938 185210 475174
rect 185446 474938 215930 475174
rect 216166 474938 246650 475174
rect 246886 474938 277370 475174
rect 277606 474938 308090 475174
rect 308326 474938 338810 475174
rect 339046 474938 369530 475174
rect 369766 474938 400250 475174
rect 400486 474938 430970 475174
rect 431206 474938 461690 475174
rect 461926 474938 492410 475174
rect 492646 474938 523130 475174
rect 523366 474938 553850 475174
rect 554086 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 586302 475174
rect 586538 474938 586622 475174
rect 586858 474938 592650 475174
rect -8726 474854 592650 474938
rect -8726 474618 -2934 474854
rect -2698 474618 -2614 474854
rect -2378 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 31610 474854
rect 31846 474618 62330 474854
rect 62566 474618 93050 474854
rect 93286 474618 123770 474854
rect 124006 474618 154490 474854
rect 154726 474618 185210 474854
rect 185446 474618 215930 474854
rect 216166 474618 246650 474854
rect 246886 474618 277370 474854
rect 277606 474618 308090 474854
rect 308326 474618 338810 474854
rect 339046 474618 369530 474854
rect 369766 474618 400250 474854
rect 400486 474618 430970 474854
rect 431206 474618 461690 474854
rect 461926 474618 492410 474854
rect 492646 474618 523130 474854
rect 523366 474618 553850 474854
rect 554086 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 586302 474854
rect 586538 474618 586622 474854
rect 586858 474618 592650 474854
rect -8726 474586 592650 474618
rect -8726 471454 592650 471486
rect -8726 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 16250 471454
rect 16486 471218 46970 471454
rect 47206 471218 77690 471454
rect 77926 471218 108410 471454
rect 108646 471218 139130 471454
rect 139366 471218 169850 471454
rect 170086 471218 200570 471454
rect 200806 471218 231290 471454
rect 231526 471218 262010 471454
rect 262246 471218 292730 471454
rect 292966 471218 323450 471454
rect 323686 471218 354170 471454
rect 354406 471218 384890 471454
rect 385126 471218 415610 471454
rect 415846 471218 446330 471454
rect 446566 471218 477050 471454
rect 477286 471218 507770 471454
rect 508006 471218 538490 471454
rect 538726 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 592650 471454
rect -8726 471134 592650 471218
rect -8726 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 16250 471134
rect 16486 470898 46970 471134
rect 47206 470898 77690 471134
rect 77926 470898 108410 471134
rect 108646 470898 139130 471134
rect 139366 470898 169850 471134
rect 170086 470898 200570 471134
rect 200806 470898 231290 471134
rect 231526 470898 262010 471134
rect 262246 470898 292730 471134
rect 292966 470898 323450 471134
rect 323686 470898 354170 471134
rect 354406 470898 384890 471134
rect 385126 470898 415610 471134
rect 415846 470898 446330 471134
rect 446566 470898 477050 471134
rect 477286 470898 507770 471134
rect 508006 470898 538490 471134
rect 538726 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 592650 471134
rect -8726 470866 592650 470898
rect -8726 461494 592650 461526
rect -8726 461258 -8694 461494
rect -8458 461258 -8374 461494
rect -8138 461258 567866 461494
rect 568102 461258 568186 461494
rect 568422 461258 592062 461494
rect 592298 461258 592382 461494
rect 592618 461258 592650 461494
rect -8726 461174 592650 461258
rect -8726 460938 -8694 461174
rect -8458 460938 -8374 461174
rect -8138 460938 567866 461174
rect 568102 460938 568186 461174
rect 568422 460938 592062 461174
rect 592298 460938 592382 461174
rect 592618 460938 592650 461174
rect -8726 460906 592650 460938
rect -8726 457774 592650 457806
rect -8726 457538 -7734 457774
rect -7498 457538 -7414 457774
rect -7178 457538 591102 457774
rect 591338 457538 591422 457774
rect 591658 457538 592650 457774
rect -8726 457454 592650 457538
rect -8726 457218 -7734 457454
rect -7498 457218 -7414 457454
rect -7178 457218 591102 457454
rect 591338 457218 591422 457454
rect 591658 457218 592650 457454
rect -8726 457186 592650 457218
rect -8726 454054 592650 454086
rect -8726 453818 -6774 454054
rect -6538 453818 -6454 454054
rect -6218 453818 590142 454054
rect 590378 453818 590462 454054
rect 590698 453818 592650 454054
rect -8726 453734 592650 453818
rect -8726 453498 -6774 453734
rect -6538 453498 -6454 453734
rect -6218 453498 590142 453734
rect 590378 453498 590462 453734
rect 590698 453498 592650 453734
rect -8726 453466 592650 453498
rect -8726 450334 592650 450366
rect -8726 450098 -5814 450334
rect -5578 450098 -5494 450334
rect -5258 450098 589182 450334
rect 589418 450098 589502 450334
rect 589738 450098 592650 450334
rect -8726 450014 592650 450098
rect -8726 449778 -5814 450014
rect -5578 449778 -5494 450014
rect -5258 449778 589182 450014
rect 589418 449778 589502 450014
rect 589738 449778 592650 450014
rect -8726 449746 592650 449778
rect -8726 446614 592650 446646
rect -8726 446378 -4854 446614
rect -4618 446378 -4534 446614
rect -4298 446378 588222 446614
rect 588458 446378 588542 446614
rect 588778 446378 592650 446614
rect -8726 446294 592650 446378
rect -8726 446058 -4854 446294
rect -4618 446058 -4534 446294
rect -4298 446058 588222 446294
rect 588458 446058 588542 446294
rect 588778 446058 592650 446294
rect -8726 446026 592650 446058
rect -8726 442894 592650 442926
rect -8726 442658 -3894 442894
rect -3658 442658 -3574 442894
rect -3338 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 587262 442894
rect 587498 442658 587582 442894
rect 587818 442658 592650 442894
rect -8726 442574 592650 442658
rect -8726 442338 -3894 442574
rect -3658 442338 -3574 442574
rect -3338 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 587262 442574
rect 587498 442338 587582 442574
rect 587818 442338 592650 442574
rect -8726 442306 592650 442338
rect -8726 439174 592650 439206
rect -8726 438938 -2934 439174
rect -2698 438938 -2614 439174
rect -2378 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 31610 439174
rect 31846 438938 62330 439174
rect 62566 438938 93050 439174
rect 93286 438938 123770 439174
rect 124006 438938 154490 439174
rect 154726 438938 185210 439174
rect 185446 438938 215930 439174
rect 216166 438938 246650 439174
rect 246886 438938 277370 439174
rect 277606 438938 308090 439174
rect 308326 438938 338810 439174
rect 339046 438938 369530 439174
rect 369766 438938 400250 439174
rect 400486 438938 430970 439174
rect 431206 438938 461690 439174
rect 461926 438938 492410 439174
rect 492646 438938 523130 439174
rect 523366 438938 553850 439174
rect 554086 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 586302 439174
rect 586538 438938 586622 439174
rect 586858 438938 592650 439174
rect -8726 438854 592650 438938
rect -8726 438618 -2934 438854
rect -2698 438618 -2614 438854
rect -2378 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 31610 438854
rect 31846 438618 62330 438854
rect 62566 438618 93050 438854
rect 93286 438618 123770 438854
rect 124006 438618 154490 438854
rect 154726 438618 185210 438854
rect 185446 438618 215930 438854
rect 216166 438618 246650 438854
rect 246886 438618 277370 438854
rect 277606 438618 308090 438854
rect 308326 438618 338810 438854
rect 339046 438618 369530 438854
rect 369766 438618 400250 438854
rect 400486 438618 430970 438854
rect 431206 438618 461690 438854
rect 461926 438618 492410 438854
rect 492646 438618 523130 438854
rect 523366 438618 553850 438854
rect 554086 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 586302 438854
rect 586538 438618 586622 438854
rect 586858 438618 592650 438854
rect -8726 438586 592650 438618
rect -8726 435454 592650 435486
rect -8726 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 16250 435454
rect 16486 435218 46970 435454
rect 47206 435218 77690 435454
rect 77926 435218 108410 435454
rect 108646 435218 139130 435454
rect 139366 435218 169850 435454
rect 170086 435218 200570 435454
rect 200806 435218 231290 435454
rect 231526 435218 262010 435454
rect 262246 435218 292730 435454
rect 292966 435218 323450 435454
rect 323686 435218 354170 435454
rect 354406 435218 384890 435454
rect 385126 435218 415610 435454
rect 415846 435218 446330 435454
rect 446566 435218 477050 435454
rect 477286 435218 507770 435454
rect 508006 435218 538490 435454
rect 538726 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 592650 435454
rect -8726 435134 592650 435218
rect -8726 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 16250 435134
rect 16486 434898 46970 435134
rect 47206 434898 77690 435134
rect 77926 434898 108410 435134
rect 108646 434898 139130 435134
rect 139366 434898 169850 435134
rect 170086 434898 200570 435134
rect 200806 434898 231290 435134
rect 231526 434898 262010 435134
rect 262246 434898 292730 435134
rect 292966 434898 323450 435134
rect 323686 434898 354170 435134
rect 354406 434898 384890 435134
rect 385126 434898 415610 435134
rect 415846 434898 446330 435134
rect 446566 434898 477050 435134
rect 477286 434898 507770 435134
rect 508006 434898 538490 435134
rect 538726 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 592650 435134
rect -8726 434866 592650 434898
rect -8726 425494 592650 425526
rect -8726 425258 -8694 425494
rect -8458 425258 -8374 425494
rect -8138 425258 567866 425494
rect 568102 425258 568186 425494
rect 568422 425258 592062 425494
rect 592298 425258 592382 425494
rect 592618 425258 592650 425494
rect -8726 425174 592650 425258
rect -8726 424938 -8694 425174
rect -8458 424938 -8374 425174
rect -8138 424938 567866 425174
rect 568102 424938 568186 425174
rect 568422 424938 592062 425174
rect 592298 424938 592382 425174
rect 592618 424938 592650 425174
rect -8726 424906 592650 424938
rect -8726 421774 592650 421806
rect -8726 421538 -7734 421774
rect -7498 421538 -7414 421774
rect -7178 421538 591102 421774
rect 591338 421538 591422 421774
rect 591658 421538 592650 421774
rect -8726 421454 592650 421538
rect -8726 421218 -7734 421454
rect -7498 421218 -7414 421454
rect -7178 421218 591102 421454
rect 591338 421218 591422 421454
rect 591658 421218 592650 421454
rect -8726 421186 592650 421218
rect -8726 418054 592650 418086
rect -8726 417818 -6774 418054
rect -6538 417818 -6454 418054
rect -6218 417818 590142 418054
rect 590378 417818 590462 418054
rect 590698 417818 592650 418054
rect -8726 417734 592650 417818
rect -8726 417498 -6774 417734
rect -6538 417498 -6454 417734
rect -6218 417498 590142 417734
rect 590378 417498 590462 417734
rect 590698 417498 592650 417734
rect -8726 417466 592650 417498
rect -8726 414334 592650 414366
rect -8726 414098 -5814 414334
rect -5578 414098 -5494 414334
rect -5258 414098 589182 414334
rect 589418 414098 589502 414334
rect 589738 414098 592650 414334
rect -8726 414014 592650 414098
rect -8726 413778 -5814 414014
rect -5578 413778 -5494 414014
rect -5258 413778 589182 414014
rect 589418 413778 589502 414014
rect 589738 413778 592650 414014
rect -8726 413746 592650 413778
rect -8726 410614 592650 410646
rect -8726 410378 -4854 410614
rect -4618 410378 -4534 410614
rect -4298 410378 588222 410614
rect 588458 410378 588542 410614
rect 588778 410378 592650 410614
rect -8726 410294 592650 410378
rect -8726 410058 -4854 410294
rect -4618 410058 -4534 410294
rect -4298 410058 588222 410294
rect 588458 410058 588542 410294
rect 588778 410058 592650 410294
rect -8726 410026 592650 410058
rect -8726 406894 592650 406926
rect -8726 406658 -3894 406894
rect -3658 406658 -3574 406894
rect -3338 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 587262 406894
rect 587498 406658 587582 406894
rect 587818 406658 592650 406894
rect -8726 406574 592650 406658
rect -8726 406338 -3894 406574
rect -3658 406338 -3574 406574
rect -3338 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 587262 406574
rect 587498 406338 587582 406574
rect 587818 406338 592650 406574
rect -8726 406306 592650 406338
rect -8726 403174 592650 403206
rect -8726 402938 -2934 403174
rect -2698 402938 -2614 403174
rect -2378 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 31610 403174
rect 31846 402938 62330 403174
rect 62566 402938 93050 403174
rect 93286 402938 123770 403174
rect 124006 402938 154490 403174
rect 154726 402938 185210 403174
rect 185446 402938 215930 403174
rect 216166 402938 246650 403174
rect 246886 402938 277370 403174
rect 277606 402938 308090 403174
rect 308326 402938 338810 403174
rect 339046 402938 369530 403174
rect 369766 402938 400250 403174
rect 400486 402938 430970 403174
rect 431206 402938 461690 403174
rect 461926 402938 492410 403174
rect 492646 402938 523130 403174
rect 523366 402938 553850 403174
rect 554086 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 586302 403174
rect 586538 402938 586622 403174
rect 586858 402938 592650 403174
rect -8726 402854 592650 402938
rect -8726 402618 -2934 402854
rect -2698 402618 -2614 402854
rect -2378 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 31610 402854
rect 31846 402618 62330 402854
rect 62566 402618 93050 402854
rect 93286 402618 123770 402854
rect 124006 402618 154490 402854
rect 154726 402618 185210 402854
rect 185446 402618 215930 402854
rect 216166 402618 246650 402854
rect 246886 402618 277370 402854
rect 277606 402618 308090 402854
rect 308326 402618 338810 402854
rect 339046 402618 369530 402854
rect 369766 402618 400250 402854
rect 400486 402618 430970 402854
rect 431206 402618 461690 402854
rect 461926 402618 492410 402854
rect 492646 402618 523130 402854
rect 523366 402618 553850 402854
rect 554086 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 586302 402854
rect 586538 402618 586622 402854
rect 586858 402618 592650 402854
rect -8726 402586 592650 402618
rect -8726 399454 592650 399486
rect -8726 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 16250 399454
rect 16486 399218 46970 399454
rect 47206 399218 77690 399454
rect 77926 399218 108410 399454
rect 108646 399218 139130 399454
rect 139366 399218 169850 399454
rect 170086 399218 200570 399454
rect 200806 399218 231290 399454
rect 231526 399218 262010 399454
rect 262246 399218 292730 399454
rect 292966 399218 323450 399454
rect 323686 399218 354170 399454
rect 354406 399218 384890 399454
rect 385126 399218 415610 399454
rect 415846 399218 446330 399454
rect 446566 399218 477050 399454
rect 477286 399218 507770 399454
rect 508006 399218 538490 399454
rect 538726 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 592650 399454
rect -8726 399134 592650 399218
rect -8726 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 16250 399134
rect 16486 398898 46970 399134
rect 47206 398898 77690 399134
rect 77926 398898 108410 399134
rect 108646 398898 139130 399134
rect 139366 398898 169850 399134
rect 170086 398898 200570 399134
rect 200806 398898 231290 399134
rect 231526 398898 262010 399134
rect 262246 398898 292730 399134
rect 292966 398898 323450 399134
rect 323686 398898 354170 399134
rect 354406 398898 384890 399134
rect 385126 398898 415610 399134
rect 415846 398898 446330 399134
rect 446566 398898 477050 399134
rect 477286 398898 507770 399134
rect 508006 398898 538490 399134
rect 538726 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 592650 399134
rect -8726 398866 592650 398898
rect -8726 389494 592650 389526
rect -8726 389258 -8694 389494
rect -8458 389258 -8374 389494
rect -8138 389258 567866 389494
rect 568102 389258 568186 389494
rect 568422 389258 592062 389494
rect 592298 389258 592382 389494
rect 592618 389258 592650 389494
rect -8726 389174 592650 389258
rect -8726 388938 -8694 389174
rect -8458 388938 -8374 389174
rect -8138 388938 567866 389174
rect 568102 388938 568186 389174
rect 568422 388938 592062 389174
rect 592298 388938 592382 389174
rect 592618 388938 592650 389174
rect -8726 388906 592650 388938
rect -8726 385774 592650 385806
rect -8726 385538 -7734 385774
rect -7498 385538 -7414 385774
rect -7178 385538 591102 385774
rect 591338 385538 591422 385774
rect 591658 385538 592650 385774
rect -8726 385454 592650 385538
rect -8726 385218 -7734 385454
rect -7498 385218 -7414 385454
rect -7178 385218 591102 385454
rect 591338 385218 591422 385454
rect 591658 385218 592650 385454
rect -8726 385186 592650 385218
rect -8726 382054 592650 382086
rect -8726 381818 -6774 382054
rect -6538 381818 -6454 382054
rect -6218 381818 590142 382054
rect 590378 381818 590462 382054
rect 590698 381818 592650 382054
rect -8726 381734 592650 381818
rect -8726 381498 -6774 381734
rect -6538 381498 -6454 381734
rect -6218 381498 590142 381734
rect 590378 381498 590462 381734
rect 590698 381498 592650 381734
rect -8726 381466 592650 381498
rect -8726 378334 592650 378366
rect -8726 378098 -5814 378334
rect -5578 378098 -5494 378334
rect -5258 378098 589182 378334
rect 589418 378098 589502 378334
rect 589738 378098 592650 378334
rect -8726 378014 592650 378098
rect -8726 377778 -5814 378014
rect -5578 377778 -5494 378014
rect -5258 377778 589182 378014
rect 589418 377778 589502 378014
rect 589738 377778 592650 378014
rect -8726 377746 592650 377778
rect -8726 374614 592650 374646
rect -8726 374378 -4854 374614
rect -4618 374378 -4534 374614
rect -4298 374378 588222 374614
rect 588458 374378 588542 374614
rect 588778 374378 592650 374614
rect -8726 374294 592650 374378
rect -8726 374058 -4854 374294
rect -4618 374058 -4534 374294
rect -4298 374058 588222 374294
rect 588458 374058 588542 374294
rect 588778 374058 592650 374294
rect -8726 374026 592650 374058
rect -8726 370894 592650 370926
rect -8726 370658 -3894 370894
rect -3658 370658 -3574 370894
rect -3338 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 587262 370894
rect 587498 370658 587582 370894
rect 587818 370658 592650 370894
rect -8726 370574 592650 370658
rect -8726 370338 -3894 370574
rect -3658 370338 -3574 370574
rect -3338 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 587262 370574
rect 587498 370338 587582 370574
rect 587818 370338 592650 370574
rect -8726 370306 592650 370338
rect -8726 367174 592650 367206
rect -8726 366938 -2934 367174
rect -2698 366938 -2614 367174
rect -2378 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 31610 367174
rect 31846 366938 62330 367174
rect 62566 366938 93050 367174
rect 93286 366938 123770 367174
rect 124006 366938 154490 367174
rect 154726 366938 185210 367174
rect 185446 366938 215930 367174
rect 216166 366938 246650 367174
rect 246886 366938 277370 367174
rect 277606 366938 308090 367174
rect 308326 366938 338810 367174
rect 339046 366938 369530 367174
rect 369766 366938 400250 367174
rect 400486 366938 430970 367174
rect 431206 366938 461690 367174
rect 461926 366938 492410 367174
rect 492646 366938 523130 367174
rect 523366 366938 553850 367174
rect 554086 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 586302 367174
rect 586538 366938 586622 367174
rect 586858 366938 592650 367174
rect -8726 366854 592650 366938
rect -8726 366618 -2934 366854
rect -2698 366618 -2614 366854
rect -2378 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 31610 366854
rect 31846 366618 62330 366854
rect 62566 366618 93050 366854
rect 93286 366618 123770 366854
rect 124006 366618 154490 366854
rect 154726 366618 185210 366854
rect 185446 366618 215930 366854
rect 216166 366618 246650 366854
rect 246886 366618 277370 366854
rect 277606 366618 308090 366854
rect 308326 366618 338810 366854
rect 339046 366618 369530 366854
rect 369766 366618 400250 366854
rect 400486 366618 430970 366854
rect 431206 366618 461690 366854
rect 461926 366618 492410 366854
rect 492646 366618 523130 366854
rect 523366 366618 553850 366854
rect 554086 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 586302 366854
rect 586538 366618 586622 366854
rect 586858 366618 592650 366854
rect -8726 366586 592650 366618
rect -8726 363454 592650 363486
rect -8726 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 16250 363454
rect 16486 363218 46970 363454
rect 47206 363218 77690 363454
rect 77926 363218 108410 363454
rect 108646 363218 139130 363454
rect 139366 363218 169850 363454
rect 170086 363218 200570 363454
rect 200806 363218 231290 363454
rect 231526 363218 262010 363454
rect 262246 363218 292730 363454
rect 292966 363218 323450 363454
rect 323686 363218 354170 363454
rect 354406 363218 384890 363454
rect 385126 363218 415610 363454
rect 415846 363218 446330 363454
rect 446566 363218 477050 363454
rect 477286 363218 507770 363454
rect 508006 363218 538490 363454
rect 538726 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 592650 363454
rect -8726 363134 592650 363218
rect -8726 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 16250 363134
rect 16486 362898 46970 363134
rect 47206 362898 77690 363134
rect 77926 362898 108410 363134
rect 108646 362898 139130 363134
rect 139366 362898 169850 363134
rect 170086 362898 200570 363134
rect 200806 362898 231290 363134
rect 231526 362898 262010 363134
rect 262246 362898 292730 363134
rect 292966 362898 323450 363134
rect 323686 362898 354170 363134
rect 354406 362898 384890 363134
rect 385126 362898 415610 363134
rect 415846 362898 446330 363134
rect 446566 362898 477050 363134
rect 477286 362898 507770 363134
rect 508006 362898 538490 363134
rect 538726 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 592650 363134
rect -8726 362866 592650 362898
rect -8726 353494 592650 353526
rect -8726 353258 -8694 353494
rect -8458 353258 -8374 353494
rect -8138 353258 567866 353494
rect 568102 353258 568186 353494
rect 568422 353258 592062 353494
rect 592298 353258 592382 353494
rect 592618 353258 592650 353494
rect -8726 353174 592650 353258
rect -8726 352938 -8694 353174
rect -8458 352938 -8374 353174
rect -8138 352938 567866 353174
rect 568102 352938 568186 353174
rect 568422 352938 592062 353174
rect 592298 352938 592382 353174
rect 592618 352938 592650 353174
rect -8726 352906 592650 352938
rect -8726 349774 592650 349806
rect -8726 349538 -7734 349774
rect -7498 349538 -7414 349774
rect -7178 349538 591102 349774
rect 591338 349538 591422 349774
rect 591658 349538 592650 349774
rect -8726 349454 592650 349538
rect -8726 349218 -7734 349454
rect -7498 349218 -7414 349454
rect -7178 349218 591102 349454
rect 591338 349218 591422 349454
rect 591658 349218 592650 349454
rect -8726 349186 592650 349218
rect -8726 346054 592650 346086
rect -8726 345818 -6774 346054
rect -6538 345818 -6454 346054
rect -6218 345818 590142 346054
rect 590378 345818 590462 346054
rect 590698 345818 592650 346054
rect -8726 345734 592650 345818
rect -8726 345498 -6774 345734
rect -6538 345498 -6454 345734
rect -6218 345498 590142 345734
rect 590378 345498 590462 345734
rect 590698 345498 592650 345734
rect -8726 345466 592650 345498
rect -8726 342334 592650 342366
rect -8726 342098 -5814 342334
rect -5578 342098 -5494 342334
rect -5258 342098 589182 342334
rect 589418 342098 589502 342334
rect 589738 342098 592650 342334
rect -8726 342014 592650 342098
rect -8726 341778 -5814 342014
rect -5578 341778 -5494 342014
rect -5258 341778 589182 342014
rect 589418 341778 589502 342014
rect 589738 341778 592650 342014
rect -8726 341746 592650 341778
rect -8726 338614 592650 338646
rect -8726 338378 -4854 338614
rect -4618 338378 -4534 338614
rect -4298 338378 588222 338614
rect 588458 338378 588542 338614
rect 588778 338378 592650 338614
rect -8726 338294 592650 338378
rect -8726 338058 -4854 338294
rect -4618 338058 -4534 338294
rect -4298 338058 588222 338294
rect 588458 338058 588542 338294
rect 588778 338058 592650 338294
rect -8726 338026 592650 338058
rect -8726 334894 592650 334926
rect -8726 334658 -3894 334894
rect -3658 334658 -3574 334894
rect -3338 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 587262 334894
rect 587498 334658 587582 334894
rect 587818 334658 592650 334894
rect -8726 334574 592650 334658
rect -8726 334338 -3894 334574
rect -3658 334338 -3574 334574
rect -3338 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 587262 334574
rect 587498 334338 587582 334574
rect 587818 334338 592650 334574
rect -8726 334306 592650 334338
rect -8726 331174 592650 331206
rect -8726 330938 -2934 331174
rect -2698 330938 -2614 331174
rect -2378 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 31610 331174
rect 31846 330938 62330 331174
rect 62566 330938 93050 331174
rect 93286 330938 123770 331174
rect 124006 330938 154490 331174
rect 154726 330938 185210 331174
rect 185446 330938 215930 331174
rect 216166 330938 246650 331174
rect 246886 330938 277370 331174
rect 277606 330938 308090 331174
rect 308326 330938 338810 331174
rect 339046 330938 369530 331174
rect 369766 330938 400250 331174
rect 400486 330938 430970 331174
rect 431206 330938 461690 331174
rect 461926 330938 492410 331174
rect 492646 330938 523130 331174
rect 523366 330938 553850 331174
rect 554086 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 586302 331174
rect 586538 330938 586622 331174
rect 586858 330938 592650 331174
rect -8726 330854 592650 330938
rect -8726 330618 -2934 330854
rect -2698 330618 -2614 330854
rect -2378 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 31610 330854
rect 31846 330618 62330 330854
rect 62566 330618 93050 330854
rect 93286 330618 123770 330854
rect 124006 330618 154490 330854
rect 154726 330618 185210 330854
rect 185446 330618 215930 330854
rect 216166 330618 246650 330854
rect 246886 330618 277370 330854
rect 277606 330618 308090 330854
rect 308326 330618 338810 330854
rect 339046 330618 369530 330854
rect 369766 330618 400250 330854
rect 400486 330618 430970 330854
rect 431206 330618 461690 330854
rect 461926 330618 492410 330854
rect 492646 330618 523130 330854
rect 523366 330618 553850 330854
rect 554086 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 586302 330854
rect 586538 330618 586622 330854
rect 586858 330618 592650 330854
rect -8726 330586 592650 330618
rect -8726 327454 592650 327486
rect -8726 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 16250 327454
rect 16486 327218 46970 327454
rect 47206 327218 77690 327454
rect 77926 327218 108410 327454
rect 108646 327218 139130 327454
rect 139366 327218 169850 327454
rect 170086 327218 200570 327454
rect 200806 327218 231290 327454
rect 231526 327218 262010 327454
rect 262246 327218 292730 327454
rect 292966 327218 323450 327454
rect 323686 327218 354170 327454
rect 354406 327218 384890 327454
rect 385126 327218 415610 327454
rect 415846 327218 446330 327454
rect 446566 327218 477050 327454
rect 477286 327218 507770 327454
rect 508006 327218 538490 327454
rect 538726 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 592650 327454
rect -8726 327134 592650 327218
rect -8726 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 16250 327134
rect 16486 326898 46970 327134
rect 47206 326898 77690 327134
rect 77926 326898 108410 327134
rect 108646 326898 139130 327134
rect 139366 326898 169850 327134
rect 170086 326898 200570 327134
rect 200806 326898 231290 327134
rect 231526 326898 262010 327134
rect 262246 326898 292730 327134
rect 292966 326898 323450 327134
rect 323686 326898 354170 327134
rect 354406 326898 384890 327134
rect 385126 326898 415610 327134
rect 415846 326898 446330 327134
rect 446566 326898 477050 327134
rect 477286 326898 507770 327134
rect 508006 326898 538490 327134
rect 538726 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 592650 327134
rect -8726 326866 592650 326898
rect -8726 317494 592650 317526
rect -8726 317258 -8694 317494
rect -8458 317258 -8374 317494
rect -8138 317258 567866 317494
rect 568102 317258 568186 317494
rect 568422 317258 592062 317494
rect 592298 317258 592382 317494
rect 592618 317258 592650 317494
rect -8726 317174 592650 317258
rect -8726 316938 -8694 317174
rect -8458 316938 -8374 317174
rect -8138 316938 567866 317174
rect 568102 316938 568186 317174
rect 568422 316938 592062 317174
rect 592298 316938 592382 317174
rect 592618 316938 592650 317174
rect -8726 316906 592650 316938
rect -8726 313774 592650 313806
rect -8726 313538 -7734 313774
rect -7498 313538 -7414 313774
rect -7178 313538 591102 313774
rect 591338 313538 591422 313774
rect 591658 313538 592650 313774
rect -8726 313454 592650 313538
rect -8726 313218 -7734 313454
rect -7498 313218 -7414 313454
rect -7178 313218 591102 313454
rect 591338 313218 591422 313454
rect 591658 313218 592650 313454
rect -8726 313186 592650 313218
rect -8726 310054 592650 310086
rect -8726 309818 -6774 310054
rect -6538 309818 -6454 310054
rect -6218 309818 590142 310054
rect 590378 309818 590462 310054
rect 590698 309818 592650 310054
rect -8726 309734 592650 309818
rect -8726 309498 -6774 309734
rect -6538 309498 -6454 309734
rect -6218 309498 590142 309734
rect 590378 309498 590462 309734
rect 590698 309498 592650 309734
rect -8726 309466 592650 309498
rect -8726 306334 592650 306366
rect -8726 306098 -5814 306334
rect -5578 306098 -5494 306334
rect -5258 306098 589182 306334
rect 589418 306098 589502 306334
rect 589738 306098 592650 306334
rect -8726 306014 592650 306098
rect -8726 305778 -5814 306014
rect -5578 305778 -5494 306014
rect -5258 305778 589182 306014
rect 589418 305778 589502 306014
rect 589738 305778 592650 306014
rect -8726 305746 592650 305778
rect -8726 302614 592650 302646
rect -8726 302378 -4854 302614
rect -4618 302378 -4534 302614
rect -4298 302378 588222 302614
rect 588458 302378 588542 302614
rect 588778 302378 592650 302614
rect -8726 302294 592650 302378
rect -8726 302058 -4854 302294
rect -4618 302058 -4534 302294
rect -4298 302058 588222 302294
rect 588458 302058 588542 302294
rect 588778 302058 592650 302294
rect -8726 302026 592650 302058
rect -8726 298894 592650 298926
rect -8726 298658 -3894 298894
rect -3658 298658 -3574 298894
rect -3338 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 587262 298894
rect 587498 298658 587582 298894
rect 587818 298658 592650 298894
rect -8726 298574 592650 298658
rect -8726 298338 -3894 298574
rect -3658 298338 -3574 298574
rect -3338 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 587262 298574
rect 587498 298338 587582 298574
rect 587818 298338 592650 298574
rect -8726 298306 592650 298338
rect -8726 295174 592650 295206
rect -8726 294938 -2934 295174
rect -2698 294938 -2614 295174
rect -2378 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 31610 295174
rect 31846 294938 62330 295174
rect 62566 294938 93050 295174
rect 93286 294938 123770 295174
rect 124006 294938 154490 295174
rect 154726 294938 185210 295174
rect 185446 294938 215930 295174
rect 216166 294938 246650 295174
rect 246886 294938 277370 295174
rect 277606 294938 308090 295174
rect 308326 294938 338810 295174
rect 339046 294938 369530 295174
rect 369766 294938 400250 295174
rect 400486 294938 430970 295174
rect 431206 294938 461690 295174
rect 461926 294938 492410 295174
rect 492646 294938 523130 295174
rect 523366 294938 553850 295174
rect 554086 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 586302 295174
rect 586538 294938 586622 295174
rect 586858 294938 592650 295174
rect -8726 294854 592650 294938
rect -8726 294618 -2934 294854
rect -2698 294618 -2614 294854
rect -2378 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 31610 294854
rect 31846 294618 62330 294854
rect 62566 294618 93050 294854
rect 93286 294618 123770 294854
rect 124006 294618 154490 294854
rect 154726 294618 185210 294854
rect 185446 294618 215930 294854
rect 216166 294618 246650 294854
rect 246886 294618 277370 294854
rect 277606 294618 308090 294854
rect 308326 294618 338810 294854
rect 339046 294618 369530 294854
rect 369766 294618 400250 294854
rect 400486 294618 430970 294854
rect 431206 294618 461690 294854
rect 461926 294618 492410 294854
rect 492646 294618 523130 294854
rect 523366 294618 553850 294854
rect 554086 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 586302 294854
rect 586538 294618 586622 294854
rect 586858 294618 592650 294854
rect -8726 294586 592650 294618
rect -8726 291454 592650 291486
rect -8726 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 16250 291454
rect 16486 291218 46970 291454
rect 47206 291218 77690 291454
rect 77926 291218 108410 291454
rect 108646 291218 139130 291454
rect 139366 291218 169850 291454
rect 170086 291218 200570 291454
rect 200806 291218 231290 291454
rect 231526 291218 262010 291454
rect 262246 291218 292730 291454
rect 292966 291218 323450 291454
rect 323686 291218 354170 291454
rect 354406 291218 384890 291454
rect 385126 291218 415610 291454
rect 415846 291218 446330 291454
rect 446566 291218 477050 291454
rect 477286 291218 507770 291454
rect 508006 291218 538490 291454
rect 538726 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 592650 291454
rect -8726 291134 592650 291218
rect -8726 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 16250 291134
rect 16486 290898 46970 291134
rect 47206 290898 77690 291134
rect 77926 290898 108410 291134
rect 108646 290898 139130 291134
rect 139366 290898 169850 291134
rect 170086 290898 200570 291134
rect 200806 290898 231290 291134
rect 231526 290898 262010 291134
rect 262246 290898 292730 291134
rect 292966 290898 323450 291134
rect 323686 290898 354170 291134
rect 354406 290898 384890 291134
rect 385126 290898 415610 291134
rect 415846 290898 446330 291134
rect 446566 290898 477050 291134
rect 477286 290898 507770 291134
rect 508006 290898 538490 291134
rect 538726 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 592650 291134
rect -8726 290866 592650 290898
rect -8726 281494 592650 281526
rect -8726 281258 -8694 281494
rect -8458 281258 -8374 281494
rect -8138 281258 567866 281494
rect 568102 281258 568186 281494
rect 568422 281258 592062 281494
rect 592298 281258 592382 281494
rect 592618 281258 592650 281494
rect -8726 281174 592650 281258
rect -8726 280938 -8694 281174
rect -8458 280938 -8374 281174
rect -8138 280938 567866 281174
rect 568102 280938 568186 281174
rect 568422 280938 592062 281174
rect 592298 280938 592382 281174
rect 592618 280938 592650 281174
rect -8726 280906 592650 280938
rect -8726 277774 592650 277806
rect -8726 277538 -7734 277774
rect -7498 277538 -7414 277774
rect -7178 277538 591102 277774
rect 591338 277538 591422 277774
rect 591658 277538 592650 277774
rect -8726 277454 592650 277538
rect -8726 277218 -7734 277454
rect -7498 277218 -7414 277454
rect -7178 277218 591102 277454
rect 591338 277218 591422 277454
rect 591658 277218 592650 277454
rect -8726 277186 592650 277218
rect -8726 274054 592650 274086
rect -8726 273818 -6774 274054
rect -6538 273818 -6454 274054
rect -6218 273818 590142 274054
rect 590378 273818 590462 274054
rect 590698 273818 592650 274054
rect -8726 273734 592650 273818
rect -8726 273498 -6774 273734
rect -6538 273498 -6454 273734
rect -6218 273498 590142 273734
rect 590378 273498 590462 273734
rect 590698 273498 592650 273734
rect -8726 273466 592650 273498
rect -8726 270334 592650 270366
rect -8726 270098 -5814 270334
rect -5578 270098 -5494 270334
rect -5258 270098 589182 270334
rect 589418 270098 589502 270334
rect 589738 270098 592650 270334
rect -8726 270014 592650 270098
rect -8726 269778 -5814 270014
rect -5578 269778 -5494 270014
rect -5258 269778 589182 270014
rect 589418 269778 589502 270014
rect 589738 269778 592650 270014
rect -8726 269746 592650 269778
rect -8726 266614 592650 266646
rect -8726 266378 -4854 266614
rect -4618 266378 -4534 266614
rect -4298 266378 588222 266614
rect 588458 266378 588542 266614
rect 588778 266378 592650 266614
rect -8726 266294 592650 266378
rect -8726 266058 -4854 266294
rect -4618 266058 -4534 266294
rect -4298 266058 588222 266294
rect 588458 266058 588542 266294
rect 588778 266058 592650 266294
rect -8726 266026 592650 266058
rect -8726 262894 592650 262926
rect -8726 262658 -3894 262894
rect -3658 262658 -3574 262894
rect -3338 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 587262 262894
rect 587498 262658 587582 262894
rect 587818 262658 592650 262894
rect -8726 262574 592650 262658
rect -8726 262338 -3894 262574
rect -3658 262338 -3574 262574
rect -3338 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 587262 262574
rect 587498 262338 587582 262574
rect 587818 262338 592650 262574
rect -8726 262306 592650 262338
rect -8726 259174 592650 259206
rect -8726 258938 -2934 259174
rect -2698 258938 -2614 259174
rect -2378 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 31610 259174
rect 31846 258938 62330 259174
rect 62566 258938 93050 259174
rect 93286 258938 123770 259174
rect 124006 258938 154490 259174
rect 154726 258938 185210 259174
rect 185446 258938 215930 259174
rect 216166 258938 246650 259174
rect 246886 258938 277370 259174
rect 277606 258938 308090 259174
rect 308326 258938 338810 259174
rect 339046 258938 369530 259174
rect 369766 258938 400250 259174
rect 400486 258938 430970 259174
rect 431206 258938 461690 259174
rect 461926 258938 492410 259174
rect 492646 258938 523130 259174
rect 523366 258938 553850 259174
rect 554086 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 586302 259174
rect 586538 258938 586622 259174
rect 586858 258938 592650 259174
rect -8726 258854 592650 258938
rect -8726 258618 -2934 258854
rect -2698 258618 -2614 258854
rect -2378 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 31610 258854
rect 31846 258618 62330 258854
rect 62566 258618 93050 258854
rect 93286 258618 123770 258854
rect 124006 258618 154490 258854
rect 154726 258618 185210 258854
rect 185446 258618 215930 258854
rect 216166 258618 246650 258854
rect 246886 258618 277370 258854
rect 277606 258618 308090 258854
rect 308326 258618 338810 258854
rect 339046 258618 369530 258854
rect 369766 258618 400250 258854
rect 400486 258618 430970 258854
rect 431206 258618 461690 258854
rect 461926 258618 492410 258854
rect 492646 258618 523130 258854
rect 523366 258618 553850 258854
rect 554086 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 586302 258854
rect 586538 258618 586622 258854
rect 586858 258618 592650 258854
rect -8726 258586 592650 258618
rect -8726 255454 592650 255486
rect -8726 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 16250 255454
rect 16486 255218 46970 255454
rect 47206 255218 77690 255454
rect 77926 255218 108410 255454
rect 108646 255218 139130 255454
rect 139366 255218 169850 255454
rect 170086 255218 200570 255454
rect 200806 255218 231290 255454
rect 231526 255218 262010 255454
rect 262246 255218 292730 255454
rect 292966 255218 323450 255454
rect 323686 255218 354170 255454
rect 354406 255218 384890 255454
rect 385126 255218 415610 255454
rect 415846 255218 446330 255454
rect 446566 255218 477050 255454
rect 477286 255218 507770 255454
rect 508006 255218 538490 255454
rect 538726 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 592650 255454
rect -8726 255134 592650 255218
rect -8726 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 16250 255134
rect 16486 254898 46970 255134
rect 47206 254898 77690 255134
rect 77926 254898 108410 255134
rect 108646 254898 139130 255134
rect 139366 254898 169850 255134
rect 170086 254898 200570 255134
rect 200806 254898 231290 255134
rect 231526 254898 262010 255134
rect 262246 254898 292730 255134
rect 292966 254898 323450 255134
rect 323686 254898 354170 255134
rect 354406 254898 384890 255134
rect 385126 254898 415610 255134
rect 415846 254898 446330 255134
rect 446566 254898 477050 255134
rect 477286 254898 507770 255134
rect 508006 254898 538490 255134
rect 538726 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 592650 255134
rect -8726 254866 592650 254898
rect -8726 245494 592650 245526
rect -8726 245258 -8694 245494
rect -8458 245258 -8374 245494
rect -8138 245258 567866 245494
rect 568102 245258 568186 245494
rect 568422 245258 592062 245494
rect 592298 245258 592382 245494
rect 592618 245258 592650 245494
rect -8726 245174 592650 245258
rect -8726 244938 -8694 245174
rect -8458 244938 -8374 245174
rect -8138 244938 567866 245174
rect 568102 244938 568186 245174
rect 568422 244938 592062 245174
rect 592298 244938 592382 245174
rect 592618 244938 592650 245174
rect -8726 244906 592650 244938
rect -8726 241774 592650 241806
rect -8726 241538 -7734 241774
rect -7498 241538 -7414 241774
rect -7178 241538 591102 241774
rect 591338 241538 591422 241774
rect 591658 241538 592650 241774
rect -8726 241454 592650 241538
rect -8726 241218 -7734 241454
rect -7498 241218 -7414 241454
rect -7178 241218 591102 241454
rect 591338 241218 591422 241454
rect 591658 241218 592650 241454
rect -8726 241186 592650 241218
rect -8726 238054 592650 238086
rect -8726 237818 -6774 238054
rect -6538 237818 -6454 238054
rect -6218 237818 590142 238054
rect 590378 237818 590462 238054
rect 590698 237818 592650 238054
rect -8726 237734 592650 237818
rect -8726 237498 -6774 237734
rect -6538 237498 -6454 237734
rect -6218 237498 590142 237734
rect 590378 237498 590462 237734
rect 590698 237498 592650 237734
rect -8726 237466 592650 237498
rect -8726 234334 592650 234366
rect -8726 234098 -5814 234334
rect -5578 234098 -5494 234334
rect -5258 234098 589182 234334
rect 589418 234098 589502 234334
rect 589738 234098 592650 234334
rect -8726 234014 592650 234098
rect -8726 233778 -5814 234014
rect -5578 233778 -5494 234014
rect -5258 233778 589182 234014
rect 589418 233778 589502 234014
rect 589738 233778 592650 234014
rect -8726 233746 592650 233778
rect -8726 230614 592650 230646
rect -8726 230378 -4854 230614
rect -4618 230378 -4534 230614
rect -4298 230378 588222 230614
rect 588458 230378 588542 230614
rect 588778 230378 592650 230614
rect -8726 230294 592650 230378
rect -8726 230058 -4854 230294
rect -4618 230058 -4534 230294
rect -4298 230058 588222 230294
rect 588458 230058 588542 230294
rect 588778 230058 592650 230294
rect -8726 230026 592650 230058
rect -8726 226894 592650 226926
rect -8726 226658 -3894 226894
rect -3658 226658 -3574 226894
rect -3338 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 587262 226894
rect 587498 226658 587582 226894
rect 587818 226658 592650 226894
rect -8726 226574 592650 226658
rect -8726 226338 -3894 226574
rect -3658 226338 -3574 226574
rect -3338 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 587262 226574
rect 587498 226338 587582 226574
rect 587818 226338 592650 226574
rect -8726 226306 592650 226338
rect -8726 223174 592650 223206
rect -8726 222938 -2934 223174
rect -2698 222938 -2614 223174
rect -2378 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 31610 223174
rect 31846 222938 62330 223174
rect 62566 222938 93050 223174
rect 93286 222938 123770 223174
rect 124006 222938 154490 223174
rect 154726 222938 185210 223174
rect 185446 222938 215930 223174
rect 216166 222938 246650 223174
rect 246886 222938 277370 223174
rect 277606 222938 308090 223174
rect 308326 222938 338810 223174
rect 339046 222938 369530 223174
rect 369766 222938 400250 223174
rect 400486 222938 430970 223174
rect 431206 222938 461690 223174
rect 461926 222938 492410 223174
rect 492646 222938 523130 223174
rect 523366 222938 553850 223174
rect 554086 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 586302 223174
rect 586538 222938 586622 223174
rect 586858 222938 592650 223174
rect -8726 222854 592650 222938
rect -8726 222618 -2934 222854
rect -2698 222618 -2614 222854
rect -2378 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 31610 222854
rect 31846 222618 62330 222854
rect 62566 222618 93050 222854
rect 93286 222618 123770 222854
rect 124006 222618 154490 222854
rect 154726 222618 185210 222854
rect 185446 222618 215930 222854
rect 216166 222618 246650 222854
rect 246886 222618 277370 222854
rect 277606 222618 308090 222854
rect 308326 222618 338810 222854
rect 339046 222618 369530 222854
rect 369766 222618 400250 222854
rect 400486 222618 430970 222854
rect 431206 222618 461690 222854
rect 461926 222618 492410 222854
rect 492646 222618 523130 222854
rect 523366 222618 553850 222854
rect 554086 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 586302 222854
rect 586538 222618 586622 222854
rect 586858 222618 592650 222854
rect -8726 222586 592650 222618
rect -8726 219454 592650 219486
rect -8726 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 16250 219454
rect 16486 219218 46970 219454
rect 47206 219218 77690 219454
rect 77926 219218 108410 219454
rect 108646 219218 139130 219454
rect 139366 219218 169850 219454
rect 170086 219218 200570 219454
rect 200806 219218 231290 219454
rect 231526 219218 262010 219454
rect 262246 219218 292730 219454
rect 292966 219218 323450 219454
rect 323686 219218 354170 219454
rect 354406 219218 384890 219454
rect 385126 219218 415610 219454
rect 415846 219218 446330 219454
rect 446566 219218 477050 219454
rect 477286 219218 507770 219454
rect 508006 219218 538490 219454
rect 538726 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 592650 219454
rect -8726 219134 592650 219218
rect -8726 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 16250 219134
rect 16486 218898 46970 219134
rect 47206 218898 77690 219134
rect 77926 218898 108410 219134
rect 108646 218898 139130 219134
rect 139366 218898 169850 219134
rect 170086 218898 200570 219134
rect 200806 218898 231290 219134
rect 231526 218898 262010 219134
rect 262246 218898 292730 219134
rect 292966 218898 323450 219134
rect 323686 218898 354170 219134
rect 354406 218898 384890 219134
rect 385126 218898 415610 219134
rect 415846 218898 446330 219134
rect 446566 218898 477050 219134
rect 477286 218898 507770 219134
rect 508006 218898 538490 219134
rect 538726 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 592650 219134
rect -8726 218866 592650 218898
rect -8726 209494 592650 209526
rect -8726 209258 -8694 209494
rect -8458 209258 -8374 209494
rect -8138 209258 567866 209494
rect 568102 209258 568186 209494
rect 568422 209258 592062 209494
rect 592298 209258 592382 209494
rect 592618 209258 592650 209494
rect -8726 209174 592650 209258
rect -8726 208938 -8694 209174
rect -8458 208938 -8374 209174
rect -8138 208938 567866 209174
rect 568102 208938 568186 209174
rect 568422 208938 592062 209174
rect 592298 208938 592382 209174
rect 592618 208938 592650 209174
rect -8726 208906 592650 208938
rect -8726 205774 592650 205806
rect -8726 205538 -7734 205774
rect -7498 205538 -7414 205774
rect -7178 205538 591102 205774
rect 591338 205538 591422 205774
rect 591658 205538 592650 205774
rect -8726 205454 592650 205538
rect -8726 205218 -7734 205454
rect -7498 205218 -7414 205454
rect -7178 205218 591102 205454
rect 591338 205218 591422 205454
rect 591658 205218 592650 205454
rect -8726 205186 592650 205218
rect -8726 202054 592650 202086
rect -8726 201818 -6774 202054
rect -6538 201818 -6454 202054
rect -6218 201818 590142 202054
rect 590378 201818 590462 202054
rect 590698 201818 592650 202054
rect -8726 201734 592650 201818
rect -8726 201498 -6774 201734
rect -6538 201498 -6454 201734
rect -6218 201498 590142 201734
rect 590378 201498 590462 201734
rect 590698 201498 592650 201734
rect -8726 201466 592650 201498
rect -8726 198334 592650 198366
rect -8726 198098 -5814 198334
rect -5578 198098 -5494 198334
rect -5258 198098 589182 198334
rect 589418 198098 589502 198334
rect 589738 198098 592650 198334
rect -8726 198014 592650 198098
rect -8726 197778 -5814 198014
rect -5578 197778 -5494 198014
rect -5258 197778 589182 198014
rect 589418 197778 589502 198014
rect 589738 197778 592650 198014
rect -8726 197746 592650 197778
rect -8726 194614 592650 194646
rect -8726 194378 -4854 194614
rect -4618 194378 -4534 194614
rect -4298 194378 588222 194614
rect 588458 194378 588542 194614
rect 588778 194378 592650 194614
rect -8726 194294 592650 194378
rect -8726 194058 -4854 194294
rect -4618 194058 -4534 194294
rect -4298 194058 588222 194294
rect 588458 194058 588542 194294
rect 588778 194058 592650 194294
rect -8726 194026 592650 194058
rect -8726 190894 592650 190926
rect -8726 190658 -3894 190894
rect -3658 190658 -3574 190894
rect -3338 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 587262 190894
rect 587498 190658 587582 190894
rect 587818 190658 592650 190894
rect -8726 190574 592650 190658
rect -8726 190338 -3894 190574
rect -3658 190338 -3574 190574
rect -3338 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 587262 190574
rect 587498 190338 587582 190574
rect 587818 190338 592650 190574
rect -8726 190306 592650 190338
rect -8726 187174 592650 187206
rect -8726 186938 -2934 187174
rect -2698 186938 -2614 187174
rect -2378 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 31610 187174
rect 31846 186938 62330 187174
rect 62566 186938 93050 187174
rect 93286 186938 123770 187174
rect 124006 186938 154490 187174
rect 154726 186938 185210 187174
rect 185446 186938 215930 187174
rect 216166 186938 246650 187174
rect 246886 186938 277370 187174
rect 277606 186938 308090 187174
rect 308326 186938 338810 187174
rect 339046 186938 369530 187174
rect 369766 186938 400250 187174
rect 400486 186938 430970 187174
rect 431206 186938 461690 187174
rect 461926 186938 492410 187174
rect 492646 186938 523130 187174
rect 523366 186938 553850 187174
rect 554086 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 586302 187174
rect 586538 186938 586622 187174
rect 586858 186938 592650 187174
rect -8726 186854 592650 186938
rect -8726 186618 -2934 186854
rect -2698 186618 -2614 186854
rect -2378 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 31610 186854
rect 31846 186618 62330 186854
rect 62566 186618 93050 186854
rect 93286 186618 123770 186854
rect 124006 186618 154490 186854
rect 154726 186618 185210 186854
rect 185446 186618 215930 186854
rect 216166 186618 246650 186854
rect 246886 186618 277370 186854
rect 277606 186618 308090 186854
rect 308326 186618 338810 186854
rect 339046 186618 369530 186854
rect 369766 186618 400250 186854
rect 400486 186618 430970 186854
rect 431206 186618 461690 186854
rect 461926 186618 492410 186854
rect 492646 186618 523130 186854
rect 523366 186618 553850 186854
rect 554086 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 586302 186854
rect 586538 186618 586622 186854
rect 586858 186618 592650 186854
rect -8726 186586 592650 186618
rect -8726 183454 592650 183486
rect -8726 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 16250 183454
rect 16486 183218 46970 183454
rect 47206 183218 77690 183454
rect 77926 183218 108410 183454
rect 108646 183218 139130 183454
rect 139366 183218 169850 183454
rect 170086 183218 200570 183454
rect 200806 183218 231290 183454
rect 231526 183218 262010 183454
rect 262246 183218 292730 183454
rect 292966 183218 323450 183454
rect 323686 183218 354170 183454
rect 354406 183218 384890 183454
rect 385126 183218 415610 183454
rect 415846 183218 446330 183454
rect 446566 183218 477050 183454
rect 477286 183218 507770 183454
rect 508006 183218 538490 183454
rect 538726 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 592650 183454
rect -8726 183134 592650 183218
rect -8726 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 16250 183134
rect 16486 182898 46970 183134
rect 47206 182898 77690 183134
rect 77926 182898 108410 183134
rect 108646 182898 139130 183134
rect 139366 182898 169850 183134
rect 170086 182898 200570 183134
rect 200806 182898 231290 183134
rect 231526 182898 262010 183134
rect 262246 182898 292730 183134
rect 292966 182898 323450 183134
rect 323686 182898 354170 183134
rect 354406 182898 384890 183134
rect 385126 182898 415610 183134
rect 415846 182898 446330 183134
rect 446566 182898 477050 183134
rect 477286 182898 507770 183134
rect 508006 182898 538490 183134
rect 538726 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 592650 183134
rect -8726 182866 592650 182898
rect -8726 173494 592650 173526
rect -8726 173258 -8694 173494
rect -8458 173258 -8374 173494
rect -8138 173258 567866 173494
rect 568102 173258 568186 173494
rect 568422 173258 592062 173494
rect 592298 173258 592382 173494
rect 592618 173258 592650 173494
rect -8726 173174 592650 173258
rect -8726 172938 -8694 173174
rect -8458 172938 -8374 173174
rect -8138 172938 567866 173174
rect 568102 172938 568186 173174
rect 568422 172938 592062 173174
rect 592298 172938 592382 173174
rect 592618 172938 592650 173174
rect -8726 172906 592650 172938
rect -8726 169774 592650 169806
rect -8726 169538 -7734 169774
rect -7498 169538 -7414 169774
rect -7178 169538 591102 169774
rect 591338 169538 591422 169774
rect 591658 169538 592650 169774
rect -8726 169454 592650 169538
rect -8726 169218 -7734 169454
rect -7498 169218 -7414 169454
rect -7178 169218 591102 169454
rect 591338 169218 591422 169454
rect 591658 169218 592650 169454
rect -8726 169186 592650 169218
rect -8726 166054 592650 166086
rect -8726 165818 -6774 166054
rect -6538 165818 -6454 166054
rect -6218 165818 590142 166054
rect 590378 165818 590462 166054
rect 590698 165818 592650 166054
rect -8726 165734 592650 165818
rect -8726 165498 -6774 165734
rect -6538 165498 -6454 165734
rect -6218 165498 590142 165734
rect 590378 165498 590462 165734
rect 590698 165498 592650 165734
rect -8726 165466 592650 165498
rect -8726 162334 592650 162366
rect -8726 162098 -5814 162334
rect -5578 162098 -5494 162334
rect -5258 162098 589182 162334
rect 589418 162098 589502 162334
rect 589738 162098 592650 162334
rect -8726 162014 592650 162098
rect -8726 161778 -5814 162014
rect -5578 161778 -5494 162014
rect -5258 161778 589182 162014
rect 589418 161778 589502 162014
rect 589738 161778 592650 162014
rect -8726 161746 592650 161778
rect -8726 158614 592650 158646
rect -8726 158378 -4854 158614
rect -4618 158378 -4534 158614
rect -4298 158378 588222 158614
rect 588458 158378 588542 158614
rect 588778 158378 592650 158614
rect -8726 158294 592650 158378
rect -8726 158058 -4854 158294
rect -4618 158058 -4534 158294
rect -4298 158058 588222 158294
rect 588458 158058 588542 158294
rect 588778 158058 592650 158294
rect -8726 158026 592650 158058
rect -8726 154894 592650 154926
rect -8726 154658 -3894 154894
rect -3658 154658 -3574 154894
rect -3338 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 587262 154894
rect 587498 154658 587582 154894
rect 587818 154658 592650 154894
rect -8726 154574 592650 154658
rect -8726 154338 -3894 154574
rect -3658 154338 -3574 154574
rect -3338 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 587262 154574
rect 587498 154338 587582 154574
rect 587818 154338 592650 154574
rect -8726 154306 592650 154338
rect -8726 151174 592650 151206
rect -8726 150938 -2934 151174
rect -2698 150938 -2614 151174
rect -2378 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 31610 151174
rect 31846 150938 62330 151174
rect 62566 150938 93050 151174
rect 93286 150938 123770 151174
rect 124006 150938 154490 151174
rect 154726 150938 185210 151174
rect 185446 150938 215930 151174
rect 216166 150938 246650 151174
rect 246886 150938 277370 151174
rect 277606 150938 308090 151174
rect 308326 150938 338810 151174
rect 339046 150938 369530 151174
rect 369766 150938 400250 151174
rect 400486 150938 430970 151174
rect 431206 150938 461690 151174
rect 461926 150938 492410 151174
rect 492646 150938 523130 151174
rect 523366 150938 553850 151174
rect 554086 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 586302 151174
rect 586538 150938 586622 151174
rect 586858 150938 592650 151174
rect -8726 150854 592650 150938
rect -8726 150618 -2934 150854
rect -2698 150618 -2614 150854
rect -2378 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 31610 150854
rect 31846 150618 62330 150854
rect 62566 150618 93050 150854
rect 93286 150618 123770 150854
rect 124006 150618 154490 150854
rect 154726 150618 185210 150854
rect 185446 150618 215930 150854
rect 216166 150618 246650 150854
rect 246886 150618 277370 150854
rect 277606 150618 308090 150854
rect 308326 150618 338810 150854
rect 339046 150618 369530 150854
rect 369766 150618 400250 150854
rect 400486 150618 430970 150854
rect 431206 150618 461690 150854
rect 461926 150618 492410 150854
rect 492646 150618 523130 150854
rect 523366 150618 553850 150854
rect 554086 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 586302 150854
rect 586538 150618 586622 150854
rect 586858 150618 592650 150854
rect -8726 150586 592650 150618
rect -8726 147454 592650 147486
rect -8726 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 16250 147454
rect 16486 147218 46970 147454
rect 47206 147218 77690 147454
rect 77926 147218 108410 147454
rect 108646 147218 139130 147454
rect 139366 147218 169850 147454
rect 170086 147218 200570 147454
rect 200806 147218 231290 147454
rect 231526 147218 262010 147454
rect 262246 147218 292730 147454
rect 292966 147218 323450 147454
rect 323686 147218 354170 147454
rect 354406 147218 384890 147454
rect 385126 147218 415610 147454
rect 415846 147218 446330 147454
rect 446566 147218 477050 147454
rect 477286 147218 507770 147454
rect 508006 147218 538490 147454
rect 538726 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 592650 147454
rect -8726 147134 592650 147218
rect -8726 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 16250 147134
rect 16486 146898 46970 147134
rect 47206 146898 77690 147134
rect 77926 146898 108410 147134
rect 108646 146898 139130 147134
rect 139366 146898 169850 147134
rect 170086 146898 200570 147134
rect 200806 146898 231290 147134
rect 231526 146898 262010 147134
rect 262246 146898 292730 147134
rect 292966 146898 323450 147134
rect 323686 146898 354170 147134
rect 354406 146898 384890 147134
rect 385126 146898 415610 147134
rect 415846 146898 446330 147134
rect 446566 146898 477050 147134
rect 477286 146898 507770 147134
rect 508006 146898 538490 147134
rect 538726 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 592650 147134
rect -8726 146866 592650 146898
rect -8726 137494 592650 137526
rect -8726 137258 -8694 137494
rect -8458 137258 -8374 137494
rect -8138 137258 567866 137494
rect 568102 137258 568186 137494
rect 568422 137258 592062 137494
rect 592298 137258 592382 137494
rect 592618 137258 592650 137494
rect -8726 137174 592650 137258
rect -8726 136938 -8694 137174
rect -8458 136938 -8374 137174
rect -8138 136938 567866 137174
rect 568102 136938 568186 137174
rect 568422 136938 592062 137174
rect 592298 136938 592382 137174
rect 592618 136938 592650 137174
rect -8726 136906 592650 136938
rect -8726 133774 592650 133806
rect -8726 133538 -7734 133774
rect -7498 133538 -7414 133774
rect -7178 133538 591102 133774
rect 591338 133538 591422 133774
rect 591658 133538 592650 133774
rect -8726 133454 592650 133538
rect -8726 133218 -7734 133454
rect -7498 133218 -7414 133454
rect -7178 133218 591102 133454
rect 591338 133218 591422 133454
rect 591658 133218 592650 133454
rect -8726 133186 592650 133218
rect -8726 130054 592650 130086
rect -8726 129818 -6774 130054
rect -6538 129818 -6454 130054
rect -6218 129818 590142 130054
rect 590378 129818 590462 130054
rect 590698 129818 592650 130054
rect -8726 129734 592650 129818
rect -8726 129498 -6774 129734
rect -6538 129498 -6454 129734
rect -6218 129498 590142 129734
rect 590378 129498 590462 129734
rect 590698 129498 592650 129734
rect -8726 129466 592650 129498
rect -8726 126334 592650 126366
rect -8726 126098 -5814 126334
rect -5578 126098 -5494 126334
rect -5258 126098 589182 126334
rect 589418 126098 589502 126334
rect 589738 126098 592650 126334
rect -8726 126014 592650 126098
rect -8726 125778 -5814 126014
rect -5578 125778 -5494 126014
rect -5258 125778 589182 126014
rect 589418 125778 589502 126014
rect 589738 125778 592650 126014
rect -8726 125746 592650 125778
rect -8726 122614 592650 122646
rect -8726 122378 -4854 122614
rect -4618 122378 -4534 122614
rect -4298 122378 588222 122614
rect 588458 122378 588542 122614
rect 588778 122378 592650 122614
rect -8726 122294 592650 122378
rect -8726 122058 -4854 122294
rect -4618 122058 -4534 122294
rect -4298 122058 588222 122294
rect 588458 122058 588542 122294
rect 588778 122058 592650 122294
rect -8726 122026 592650 122058
rect -8726 118894 592650 118926
rect -8726 118658 -3894 118894
rect -3658 118658 -3574 118894
rect -3338 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 587262 118894
rect 587498 118658 587582 118894
rect 587818 118658 592650 118894
rect -8726 118574 592650 118658
rect -8726 118338 -3894 118574
rect -3658 118338 -3574 118574
rect -3338 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 587262 118574
rect 587498 118338 587582 118574
rect 587818 118338 592650 118574
rect -8726 118306 592650 118338
rect -8726 115174 592650 115206
rect -8726 114938 -2934 115174
rect -2698 114938 -2614 115174
rect -2378 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 31610 115174
rect 31846 114938 62330 115174
rect 62566 114938 93050 115174
rect 93286 114938 123770 115174
rect 124006 114938 154490 115174
rect 154726 114938 185210 115174
rect 185446 114938 215930 115174
rect 216166 114938 246650 115174
rect 246886 114938 277370 115174
rect 277606 114938 308090 115174
rect 308326 114938 338810 115174
rect 339046 114938 369530 115174
rect 369766 114938 400250 115174
rect 400486 114938 430970 115174
rect 431206 114938 461690 115174
rect 461926 114938 492410 115174
rect 492646 114938 523130 115174
rect 523366 114938 553850 115174
rect 554086 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 586302 115174
rect 586538 114938 586622 115174
rect 586858 114938 592650 115174
rect -8726 114854 592650 114938
rect -8726 114618 -2934 114854
rect -2698 114618 -2614 114854
rect -2378 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 31610 114854
rect 31846 114618 62330 114854
rect 62566 114618 93050 114854
rect 93286 114618 123770 114854
rect 124006 114618 154490 114854
rect 154726 114618 185210 114854
rect 185446 114618 215930 114854
rect 216166 114618 246650 114854
rect 246886 114618 277370 114854
rect 277606 114618 308090 114854
rect 308326 114618 338810 114854
rect 339046 114618 369530 114854
rect 369766 114618 400250 114854
rect 400486 114618 430970 114854
rect 431206 114618 461690 114854
rect 461926 114618 492410 114854
rect 492646 114618 523130 114854
rect 523366 114618 553850 114854
rect 554086 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 586302 114854
rect 586538 114618 586622 114854
rect 586858 114618 592650 114854
rect -8726 114586 592650 114618
rect -8726 111454 592650 111486
rect -8726 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 16250 111454
rect 16486 111218 46970 111454
rect 47206 111218 77690 111454
rect 77926 111218 108410 111454
rect 108646 111218 139130 111454
rect 139366 111218 169850 111454
rect 170086 111218 200570 111454
rect 200806 111218 231290 111454
rect 231526 111218 262010 111454
rect 262246 111218 292730 111454
rect 292966 111218 323450 111454
rect 323686 111218 354170 111454
rect 354406 111218 384890 111454
rect 385126 111218 415610 111454
rect 415846 111218 446330 111454
rect 446566 111218 477050 111454
rect 477286 111218 507770 111454
rect 508006 111218 538490 111454
rect 538726 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 592650 111454
rect -8726 111134 592650 111218
rect -8726 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 16250 111134
rect 16486 110898 46970 111134
rect 47206 110898 77690 111134
rect 77926 110898 108410 111134
rect 108646 110898 139130 111134
rect 139366 110898 169850 111134
rect 170086 110898 200570 111134
rect 200806 110898 231290 111134
rect 231526 110898 262010 111134
rect 262246 110898 292730 111134
rect 292966 110898 323450 111134
rect 323686 110898 354170 111134
rect 354406 110898 384890 111134
rect 385126 110898 415610 111134
rect 415846 110898 446330 111134
rect 446566 110898 477050 111134
rect 477286 110898 507770 111134
rect 508006 110898 538490 111134
rect 538726 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 592650 111134
rect -8726 110866 592650 110898
rect -8726 101494 592650 101526
rect -8726 101258 -8694 101494
rect -8458 101258 -8374 101494
rect -8138 101258 567866 101494
rect 568102 101258 568186 101494
rect 568422 101258 592062 101494
rect 592298 101258 592382 101494
rect 592618 101258 592650 101494
rect -8726 101174 592650 101258
rect -8726 100938 -8694 101174
rect -8458 100938 -8374 101174
rect -8138 100938 567866 101174
rect 568102 100938 568186 101174
rect 568422 100938 592062 101174
rect 592298 100938 592382 101174
rect 592618 100938 592650 101174
rect -8726 100906 592650 100938
rect -8726 97774 592650 97806
rect -8726 97538 -7734 97774
rect -7498 97538 -7414 97774
rect -7178 97538 591102 97774
rect 591338 97538 591422 97774
rect 591658 97538 592650 97774
rect -8726 97454 592650 97538
rect -8726 97218 -7734 97454
rect -7498 97218 -7414 97454
rect -7178 97218 591102 97454
rect 591338 97218 591422 97454
rect 591658 97218 592650 97454
rect -8726 97186 592650 97218
rect -8726 94054 592650 94086
rect -8726 93818 -6774 94054
rect -6538 93818 -6454 94054
rect -6218 93818 590142 94054
rect 590378 93818 590462 94054
rect 590698 93818 592650 94054
rect -8726 93734 592650 93818
rect -8726 93498 -6774 93734
rect -6538 93498 -6454 93734
rect -6218 93498 590142 93734
rect 590378 93498 590462 93734
rect 590698 93498 592650 93734
rect -8726 93466 592650 93498
rect -8726 90334 592650 90366
rect -8726 90098 -5814 90334
rect -5578 90098 -5494 90334
rect -5258 90098 589182 90334
rect 589418 90098 589502 90334
rect 589738 90098 592650 90334
rect -8726 90014 592650 90098
rect -8726 89778 -5814 90014
rect -5578 89778 -5494 90014
rect -5258 89778 589182 90014
rect 589418 89778 589502 90014
rect 589738 89778 592650 90014
rect -8726 89746 592650 89778
rect -8726 86614 592650 86646
rect -8726 86378 -4854 86614
rect -4618 86378 -4534 86614
rect -4298 86378 588222 86614
rect 588458 86378 588542 86614
rect 588778 86378 592650 86614
rect -8726 86294 592650 86378
rect -8726 86058 -4854 86294
rect -4618 86058 -4534 86294
rect -4298 86058 588222 86294
rect 588458 86058 588542 86294
rect 588778 86058 592650 86294
rect -8726 86026 592650 86058
rect -8726 82894 592650 82926
rect -8726 82658 -3894 82894
rect -3658 82658 -3574 82894
rect -3338 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 587262 82894
rect 587498 82658 587582 82894
rect 587818 82658 592650 82894
rect -8726 82574 592650 82658
rect -8726 82338 -3894 82574
rect -3658 82338 -3574 82574
rect -3338 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 587262 82574
rect 587498 82338 587582 82574
rect 587818 82338 592650 82574
rect -8726 82306 592650 82338
rect -8726 79174 592650 79206
rect -8726 78938 -2934 79174
rect -2698 78938 -2614 79174
rect -2378 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 31610 79174
rect 31846 78938 62330 79174
rect 62566 78938 93050 79174
rect 93286 78938 123770 79174
rect 124006 78938 154490 79174
rect 154726 78938 185210 79174
rect 185446 78938 215930 79174
rect 216166 78938 246650 79174
rect 246886 78938 277370 79174
rect 277606 78938 308090 79174
rect 308326 78938 338810 79174
rect 339046 78938 369530 79174
rect 369766 78938 400250 79174
rect 400486 78938 430970 79174
rect 431206 78938 461690 79174
rect 461926 78938 492410 79174
rect 492646 78938 523130 79174
rect 523366 78938 553850 79174
rect 554086 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 586302 79174
rect 586538 78938 586622 79174
rect 586858 78938 592650 79174
rect -8726 78854 592650 78938
rect -8726 78618 -2934 78854
rect -2698 78618 -2614 78854
rect -2378 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 31610 78854
rect 31846 78618 62330 78854
rect 62566 78618 93050 78854
rect 93286 78618 123770 78854
rect 124006 78618 154490 78854
rect 154726 78618 185210 78854
rect 185446 78618 215930 78854
rect 216166 78618 246650 78854
rect 246886 78618 277370 78854
rect 277606 78618 308090 78854
rect 308326 78618 338810 78854
rect 339046 78618 369530 78854
rect 369766 78618 400250 78854
rect 400486 78618 430970 78854
rect 431206 78618 461690 78854
rect 461926 78618 492410 78854
rect 492646 78618 523130 78854
rect 523366 78618 553850 78854
rect 554086 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 586302 78854
rect 586538 78618 586622 78854
rect 586858 78618 592650 78854
rect -8726 78586 592650 78618
rect -8726 75454 592650 75486
rect -8726 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 16250 75454
rect 16486 75218 46970 75454
rect 47206 75218 77690 75454
rect 77926 75218 108410 75454
rect 108646 75218 139130 75454
rect 139366 75218 169850 75454
rect 170086 75218 200570 75454
rect 200806 75218 231290 75454
rect 231526 75218 262010 75454
rect 262246 75218 292730 75454
rect 292966 75218 323450 75454
rect 323686 75218 354170 75454
rect 354406 75218 384890 75454
rect 385126 75218 415610 75454
rect 415846 75218 446330 75454
rect 446566 75218 477050 75454
rect 477286 75218 507770 75454
rect 508006 75218 538490 75454
rect 538726 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 592650 75454
rect -8726 75134 592650 75218
rect -8726 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 16250 75134
rect 16486 74898 46970 75134
rect 47206 74898 77690 75134
rect 77926 74898 108410 75134
rect 108646 74898 139130 75134
rect 139366 74898 169850 75134
rect 170086 74898 200570 75134
rect 200806 74898 231290 75134
rect 231526 74898 262010 75134
rect 262246 74898 292730 75134
rect 292966 74898 323450 75134
rect 323686 74898 354170 75134
rect 354406 74898 384890 75134
rect 385126 74898 415610 75134
rect 415846 74898 446330 75134
rect 446566 74898 477050 75134
rect 477286 74898 507770 75134
rect 508006 74898 538490 75134
rect 538726 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 592650 75134
rect -8726 74866 592650 74898
rect -8726 65494 592650 65526
rect -8726 65258 -8694 65494
rect -8458 65258 -8374 65494
rect -8138 65258 567866 65494
rect 568102 65258 568186 65494
rect 568422 65258 592062 65494
rect 592298 65258 592382 65494
rect 592618 65258 592650 65494
rect -8726 65174 592650 65258
rect -8726 64938 -8694 65174
rect -8458 64938 -8374 65174
rect -8138 64938 567866 65174
rect 568102 64938 568186 65174
rect 568422 64938 592062 65174
rect 592298 64938 592382 65174
rect 592618 64938 592650 65174
rect -8726 64906 592650 64938
rect -8726 61774 592650 61806
rect -8726 61538 -7734 61774
rect -7498 61538 -7414 61774
rect -7178 61538 591102 61774
rect 591338 61538 591422 61774
rect 591658 61538 592650 61774
rect -8726 61454 592650 61538
rect -8726 61218 -7734 61454
rect -7498 61218 -7414 61454
rect -7178 61218 591102 61454
rect 591338 61218 591422 61454
rect 591658 61218 592650 61454
rect -8726 61186 592650 61218
rect -8726 58054 592650 58086
rect -8726 57818 -6774 58054
rect -6538 57818 -6454 58054
rect -6218 57818 590142 58054
rect 590378 57818 590462 58054
rect 590698 57818 592650 58054
rect -8726 57734 592650 57818
rect -8726 57498 -6774 57734
rect -6538 57498 -6454 57734
rect -6218 57498 590142 57734
rect 590378 57498 590462 57734
rect 590698 57498 592650 57734
rect -8726 57466 592650 57498
rect -8726 54334 592650 54366
rect -8726 54098 -5814 54334
rect -5578 54098 -5494 54334
rect -5258 54098 589182 54334
rect 589418 54098 589502 54334
rect 589738 54098 592650 54334
rect -8726 54014 592650 54098
rect -8726 53778 -5814 54014
rect -5578 53778 -5494 54014
rect -5258 53778 589182 54014
rect 589418 53778 589502 54014
rect 589738 53778 592650 54014
rect -8726 53746 592650 53778
rect -8726 50614 592650 50646
rect -8726 50378 -4854 50614
rect -4618 50378 -4534 50614
rect -4298 50378 588222 50614
rect 588458 50378 588542 50614
rect 588778 50378 592650 50614
rect -8726 50294 592650 50378
rect -8726 50058 -4854 50294
rect -4618 50058 -4534 50294
rect -4298 50058 588222 50294
rect 588458 50058 588542 50294
rect 588778 50058 592650 50294
rect -8726 50026 592650 50058
rect -8726 46894 592650 46926
rect -8726 46658 -3894 46894
rect -3658 46658 -3574 46894
rect -3338 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 587262 46894
rect 587498 46658 587582 46894
rect 587818 46658 592650 46894
rect -8726 46574 592650 46658
rect -8726 46338 -3894 46574
rect -3658 46338 -3574 46574
rect -3338 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 587262 46574
rect 587498 46338 587582 46574
rect 587818 46338 592650 46574
rect -8726 46306 592650 46338
rect -8726 43174 592650 43206
rect -8726 42938 -2934 43174
rect -2698 42938 -2614 43174
rect -2378 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 31610 43174
rect 31846 42938 62330 43174
rect 62566 42938 93050 43174
rect 93286 42938 123770 43174
rect 124006 42938 154490 43174
rect 154726 42938 185210 43174
rect 185446 42938 215930 43174
rect 216166 42938 246650 43174
rect 246886 42938 277370 43174
rect 277606 42938 308090 43174
rect 308326 42938 338810 43174
rect 339046 42938 369530 43174
rect 369766 42938 400250 43174
rect 400486 42938 430970 43174
rect 431206 42938 461690 43174
rect 461926 42938 492410 43174
rect 492646 42938 523130 43174
rect 523366 42938 553850 43174
rect 554086 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 586302 43174
rect 586538 42938 586622 43174
rect 586858 42938 592650 43174
rect -8726 42854 592650 42938
rect -8726 42618 -2934 42854
rect -2698 42618 -2614 42854
rect -2378 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 31610 42854
rect 31846 42618 62330 42854
rect 62566 42618 93050 42854
rect 93286 42618 123770 42854
rect 124006 42618 154490 42854
rect 154726 42618 185210 42854
rect 185446 42618 215930 42854
rect 216166 42618 246650 42854
rect 246886 42618 277370 42854
rect 277606 42618 308090 42854
rect 308326 42618 338810 42854
rect 339046 42618 369530 42854
rect 369766 42618 400250 42854
rect 400486 42618 430970 42854
rect 431206 42618 461690 42854
rect 461926 42618 492410 42854
rect 492646 42618 523130 42854
rect 523366 42618 553850 42854
rect 554086 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 586302 42854
rect 586538 42618 586622 42854
rect 586858 42618 592650 42854
rect -8726 42586 592650 42618
rect -8726 39454 592650 39486
rect -8726 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 16250 39454
rect 16486 39218 46970 39454
rect 47206 39218 77690 39454
rect 77926 39218 108410 39454
rect 108646 39218 139130 39454
rect 139366 39218 169850 39454
rect 170086 39218 200570 39454
rect 200806 39218 231290 39454
rect 231526 39218 262010 39454
rect 262246 39218 292730 39454
rect 292966 39218 323450 39454
rect 323686 39218 354170 39454
rect 354406 39218 384890 39454
rect 385126 39218 415610 39454
rect 415846 39218 446330 39454
rect 446566 39218 477050 39454
rect 477286 39218 507770 39454
rect 508006 39218 538490 39454
rect 538726 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 592650 39454
rect -8726 39134 592650 39218
rect -8726 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 16250 39134
rect 16486 38898 46970 39134
rect 47206 38898 77690 39134
rect 77926 38898 108410 39134
rect 108646 38898 139130 39134
rect 139366 38898 169850 39134
rect 170086 38898 200570 39134
rect 200806 38898 231290 39134
rect 231526 38898 262010 39134
rect 262246 38898 292730 39134
rect 292966 38898 323450 39134
rect 323686 38898 354170 39134
rect 354406 38898 384890 39134
rect 385126 38898 415610 39134
rect 415846 38898 446330 39134
rect 446566 38898 477050 39134
rect 477286 38898 507770 39134
rect 508006 38898 538490 39134
rect 538726 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 592650 39134
rect -8726 38866 592650 38898
rect -8726 29494 592650 29526
rect -8726 29258 -8694 29494
rect -8458 29258 -8374 29494
rect -8138 29258 567866 29494
rect 568102 29258 568186 29494
rect 568422 29258 592062 29494
rect 592298 29258 592382 29494
rect 592618 29258 592650 29494
rect -8726 29174 592650 29258
rect -8726 28938 -8694 29174
rect -8458 28938 -8374 29174
rect -8138 28938 567866 29174
rect 568102 28938 568186 29174
rect 568422 28938 592062 29174
rect 592298 28938 592382 29174
rect 592618 28938 592650 29174
rect -8726 28906 592650 28938
rect -8726 25774 592650 25806
rect -8726 25538 -7734 25774
rect -7498 25538 -7414 25774
rect -7178 25538 591102 25774
rect 591338 25538 591422 25774
rect 591658 25538 592650 25774
rect -8726 25454 592650 25538
rect -8726 25218 -7734 25454
rect -7498 25218 -7414 25454
rect -7178 25218 591102 25454
rect 591338 25218 591422 25454
rect 591658 25218 592650 25454
rect -8726 25186 592650 25218
rect -8726 22054 592650 22086
rect -8726 21818 -6774 22054
rect -6538 21818 -6454 22054
rect -6218 21818 590142 22054
rect 590378 21818 590462 22054
rect 590698 21818 592650 22054
rect -8726 21734 592650 21818
rect -8726 21498 -6774 21734
rect -6538 21498 -6454 21734
rect -6218 21498 590142 21734
rect 590378 21498 590462 21734
rect 590698 21498 592650 21734
rect -8726 21466 592650 21498
rect -8726 18334 592650 18366
rect -8726 18098 -5814 18334
rect -5578 18098 -5494 18334
rect -5258 18098 589182 18334
rect 589418 18098 589502 18334
rect 589738 18098 592650 18334
rect -8726 18014 592650 18098
rect -8726 17778 -5814 18014
rect -5578 17778 -5494 18014
rect -5258 17778 589182 18014
rect 589418 17778 589502 18014
rect 589738 17778 592650 18014
rect -8726 17746 592650 17778
rect -8726 14614 592650 14646
rect -8726 14378 -4854 14614
rect -4618 14378 -4534 14614
rect -4298 14378 588222 14614
rect 588458 14378 588542 14614
rect 588778 14378 592650 14614
rect -8726 14294 592650 14378
rect -8726 14058 -4854 14294
rect -4618 14058 -4534 14294
rect -4298 14058 588222 14294
rect 588458 14058 588542 14294
rect 588778 14058 592650 14294
rect -8726 14026 592650 14058
rect -8726 10894 592650 10926
rect -8726 10658 -3894 10894
rect -3658 10658 -3574 10894
rect -3338 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 587262 10894
rect 587498 10658 587582 10894
rect 587818 10658 592650 10894
rect -8726 10574 592650 10658
rect -8726 10338 -3894 10574
rect -3658 10338 -3574 10574
rect -3338 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 587262 10574
rect 587498 10338 587582 10574
rect 587818 10338 592650 10574
rect -8726 10306 592650 10338
rect -8726 7174 592650 7206
rect -8726 6938 -2934 7174
rect -2698 6938 -2614 7174
rect -2378 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 586302 7174
rect 586538 6938 586622 7174
rect 586858 6938 592650 7174
rect -8726 6854 592650 6938
rect -8726 6618 -2934 6854
rect -2698 6618 -2614 6854
rect -2378 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 586302 6854
rect 586538 6618 586622 6854
rect 586858 6618 592650 6854
rect -8726 6586 592650 6618
rect -8726 3454 592650 3486
rect -8726 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 592650 3454
rect -8726 3134 592650 3218
rect -8726 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 592650 3134
rect -8726 2866 592650 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 5546 -1306
rect 5782 -1542 5866 -1306
rect 6102 -1542 41546 -1306
rect 41782 -1542 41866 -1306
rect 42102 -1542 77546 -1306
rect 77782 -1542 77866 -1306
rect 78102 -1542 113546 -1306
rect 113782 -1542 113866 -1306
rect 114102 -1542 149546 -1306
rect 149782 -1542 149866 -1306
rect 150102 -1542 185546 -1306
rect 185782 -1542 185866 -1306
rect 186102 -1542 221546 -1306
rect 221782 -1542 221866 -1306
rect 222102 -1542 257546 -1306
rect 257782 -1542 257866 -1306
rect 258102 -1542 293546 -1306
rect 293782 -1542 293866 -1306
rect 294102 -1542 329546 -1306
rect 329782 -1542 329866 -1306
rect 330102 -1542 365546 -1306
rect 365782 -1542 365866 -1306
rect 366102 -1542 401546 -1306
rect 401782 -1542 401866 -1306
rect 402102 -1542 437546 -1306
rect 437782 -1542 437866 -1306
rect 438102 -1542 473546 -1306
rect 473782 -1542 473866 -1306
rect 474102 -1542 509546 -1306
rect 509782 -1542 509866 -1306
rect 510102 -1542 545546 -1306
rect 545782 -1542 545866 -1306
rect 546102 -1542 581546 -1306
rect 581782 -1542 581866 -1306
rect 582102 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 5546 -1626
rect 5782 -1862 5866 -1626
rect 6102 -1862 41546 -1626
rect 41782 -1862 41866 -1626
rect 42102 -1862 77546 -1626
rect 77782 -1862 77866 -1626
rect 78102 -1862 113546 -1626
rect 113782 -1862 113866 -1626
rect 114102 -1862 149546 -1626
rect 149782 -1862 149866 -1626
rect 150102 -1862 185546 -1626
rect 185782 -1862 185866 -1626
rect 186102 -1862 221546 -1626
rect 221782 -1862 221866 -1626
rect 222102 -1862 257546 -1626
rect 257782 -1862 257866 -1626
rect 258102 -1862 293546 -1626
rect 293782 -1862 293866 -1626
rect 294102 -1862 329546 -1626
rect 329782 -1862 329866 -1626
rect 330102 -1862 365546 -1626
rect 365782 -1862 365866 -1626
rect 366102 -1862 401546 -1626
rect 401782 -1862 401866 -1626
rect 402102 -1862 437546 -1626
rect 437782 -1862 437866 -1626
rect 438102 -1862 473546 -1626
rect 473782 -1862 473866 -1626
rect 474102 -1862 509546 -1626
rect 509782 -1862 509866 -1626
rect 510102 -1862 545546 -1626
rect 545782 -1862 545866 -1626
rect 546102 -1862 581546 -1626
rect 581782 -1862 581866 -1626
rect 582102 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 9266 -2266
rect 9502 -2502 9586 -2266
rect 9822 -2502 45266 -2266
rect 45502 -2502 45586 -2266
rect 45822 -2502 81266 -2266
rect 81502 -2502 81586 -2266
rect 81822 -2502 117266 -2266
rect 117502 -2502 117586 -2266
rect 117822 -2502 153266 -2266
rect 153502 -2502 153586 -2266
rect 153822 -2502 189266 -2266
rect 189502 -2502 189586 -2266
rect 189822 -2502 225266 -2266
rect 225502 -2502 225586 -2266
rect 225822 -2502 261266 -2266
rect 261502 -2502 261586 -2266
rect 261822 -2502 297266 -2266
rect 297502 -2502 297586 -2266
rect 297822 -2502 333266 -2266
rect 333502 -2502 333586 -2266
rect 333822 -2502 369266 -2266
rect 369502 -2502 369586 -2266
rect 369822 -2502 405266 -2266
rect 405502 -2502 405586 -2266
rect 405822 -2502 441266 -2266
rect 441502 -2502 441586 -2266
rect 441822 -2502 477266 -2266
rect 477502 -2502 477586 -2266
rect 477822 -2502 513266 -2266
rect 513502 -2502 513586 -2266
rect 513822 -2502 549266 -2266
rect 549502 -2502 549586 -2266
rect 549822 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 9266 -2586
rect 9502 -2822 9586 -2586
rect 9822 -2822 45266 -2586
rect 45502 -2822 45586 -2586
rect 45822 -2822 81266 -2586
rect 81502 -2822 81586 -2586
rect 81822 -2822 117266 -2586
rect 117502 -2822 117586 -2586
rect 117822 -2822 153266 -2586
rect 153502 -2822 153586 -2586
rect 153822 -2822 189266 -2586
rect 189502 -2822 189586 -2586
rect 189822 -2822 225266 -2586
rect 225502 -2822 225586 -2586
rect 225822 -2822 261266 -2586
rect 261502 -2822 261586 -2586
rect 261822 -2822 297266 -2586
rect 297502 -2822 297586 -2586
rect 297822 -2822 333266 -2586
rect 333502 -2822 333586 -2586
rect 333822 -2822 369266 -2586
rect 369502 -2822 369586 -2586
rect 369822 -2822 405266 -2586
rect 405502 -2822 405586 -2586
rect 405822 -2822 441266 -2586
rect 441502 -2822 441586 -2586
rect 441822 -2822 477266 -2586
rect 477502 -2822 477586 -2586
rect 477822 -2822 513266 -2586
rect 513502 -2822 513586 -2586
rect 513822 -2822 549266 -2586
rect 549502 -2822 549586 -2586
rect 549822 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 567866 -7066
rect 568102 -7302 568186 -7066
rect 568422 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 567866 -7386
rect 568102 -7622 568186 -7386
rect 568422 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use rift2Wrap  i_Rift2Wrap
timestamp 0
transform 1 0 12000 0 1 12000
box 0 0 554204 666748
<< labels >>
flabel metal3 s 583520 285276 584960 285516 0 FreeSans 960 0 0 0 analog_io[0]
port 0 nsew signal bidirectional
flabel metal2 s 446098 703520 446210 704960 0 FreeSans 448 90 0 0 analog_io[10]
port 1 nsew signal bidirectional
flabel metal2 s 381146 703520 381258 704960 0 FreeSans 448 90 0 0 analog_io[11]
port 2 nsew signal bidirectional
flabel metal2 s 316286 703520 316398 704960 0 FreeSans 448 90 0 0 analog_io[12]
port 3 nsew signal bidirectional
flabel metal2 s 251426 703520 251538 704960 0 FreeSans 448 90 0 0 analog_io[13]
port 4 nsew signal bidirectional
flabel metal2 s 186474 703520 186586 704960 0 FreeSans 448 90 0 0 analog_io[14]
port 5 nsew signal bidirectional
flabel metal2 s 121614 703520 121726 704960 0 FreeSans 448 90 0 0 analog_io[15]
port 6 nsew signal bidirectional
flabel metal2 s 56754 703520 56866 704960 0 FreeSans 448 90 0 0 analog_io[16]
port 7 nsew signal bidirectional
flabel metal3 s -960 697220 480 697460 0 FreeSans 960 0 0 0 analog_io[17]
port 8 nsew signal bidirectional
flabel metal3 s -960 644996 480 645236 0 FreeSans 960 0 0 0 analog_io[18]
port 9 nsew signal bidirectional
flabel metal3 s -960 592908 480 593148 0 FreeSans 960 0 0 0 analog_io[19]
port 10 nsew signal bidirectional
flabel metal3 s 583520 338452 584960 338692 0 FreeSans 960 0 0 0 analog_io[1]
port 11 nsew signal bidirectional
flabel metal3 s -960 540684 480 540924 0 FreeSans 960 0 0 0 analog_io[20]
port 12 nsew signal bidirectional
flabel metal3 s -960 488596 480 488836 0 FreeSans 960 0 0 0 analog_io[21]
port 13 nsew signal bidirectional
flabel metal3 s -960 436508 480 436748 0 FreeSans 960 0 0 0 analog_io[22]
port 14 nsew signal bidirectional
flabel metal3 s -960 384284 480 384524 0 FreeSans 960 0 0 0 analog_io[23]
port 15 nsew signal bidirectional
flabel metal3 s -960 332196 480 332436 0 FreeSans 960 0 0 0 analog_io[24]
port 16 nsew signal bidirectional
flabel metal3 s -960 279972 480 280212 0 FreeSans 960 0 0 0 analog_io[25]
port 17 nsew signal bidirectional
flabel metal3 s -960 227884 480 228124 0 FreeSans 960 0 0 0 analog_io[26]
port 18 nsew signal bidirectional
flabel metal3 s -960 175796 480 176036 0 FreeSans 960 0 0 0 analog_io[27]
port 19 nsew signal bidirectional
flabel metal3 s -960 123572 480 123812 0 FreeSans 960 0 0 0 analog_io[28]
port 20 nsew signal bidirectional
flabel metal3 s 583520 391628 584960 391868 0 FreeSans 960 0 0 0 analog_io[2]
port 21 nsew signal bidirectional
flabel metal3 s 583520 444668 584960 444908 0 FreeSans 960 0 0 0 analog_io[3]
port 22 nsew signal bidirectional
flabel metal3 s 583520 497844 584960 498084 0 FreeSans 960 0 0 0 analog_io[4]
port 23 nsew signal bidirectional
flabel metal3 s 583520 551020 584960 551260 0 FreeSans 960 0 0 0 analog_io[5]
port 24 nsew signal bidirectional
flabel metal3 s 583520 604060 584960 604300 0 FreeSans 960 0 0 0 analog_io[6]
port 25 nsew signal bidirectional
flabel metal3 s 583520 657236 584960 657476 0 FreeSans 960 0 0 0 analog_io[7]
port 26 nsew signal bidirectional
flabel metal2 s 575818 703520 575930 704960 0 FreeSans 448 90 0 0 analog_io[8]
port 27 nsew signal bidirectional
flabel metal2 s 510958 703520 511070 704960 0 FreeSans 448 90 0 0 analog_io[9]
port 28 nsew signal bidirectional
flabel metal3 s 583520 6476 584960 6716 0 FreeSans 960 0 0 0 io_in[0]
port 29 nsew signal input
flabel metal3 s 583520 457996 584960 458236 0 FreeSans 960 0 0 0 io_in[10]
port 30 nsew signal input
flabel metal3 s 583520 511172 584960 511412 0 FreeSans 960 0 0 0 io_in[11]
port 31 nsew signal input
flabel metal3 s 583520 564212 584960 564452 0 FreeSans 960 0 0 0 io_in[12]
port 32 nsew signal input
flabel metal3 s 583520 617388 584960 617628 0 FreeSans 960 0 0 0 io_in[13]
port 33 nsew signal input
flabel metal3 s 583520 670564 584960 670804 0 FreeSans 960 0 0 0 io_in[14]
port 34 nsew signal input
flabel metal2 s 559626 703520 559738 704960 0 FreeSans 448 90 0 0 io_in[15]
port 35 nsew signal input
flabel metal2 s 494766 703520 494878 704960 0 FreeSans 448 90 0 0 io_in[16]
port 36 nsew signal input
flabel metal2 s 429814 703520 429926 704960 0 FreeSans 448 90 0 0 io_in[17]
port 37 nsew signal input
flabel metal2 s 364954 703520 365066 704960 0 FreeSans 448 90 0 0 io_in[18]
port 38 nsew signal input
flabel metal2 s 300094 703520 300206 704960 0 FreeSans 448 90 0 0 io_in[19]
port 39 nsew signal input
flabel metal3 s 583520 46188 584960 46428 0 FreeSans 960 0 0 0 io_in[1]
port 40 nsew signal input
flabel metal2 s 235142 703520 235254 704960 0 FreeSans 448 90 0 0 io_in[20]
port 41 nsew signal input
flabel metal2 s 170282 703520 170394 704960 0 FreeSans 448 90 0 0 io_in[21]
port 42 nsew signal input
flabel metal2 s 105422 703520 105534 704960 0 FreeSans 448 90 0 0 io_in[22]
port 43 nsew signal input
flabel metal2 s 40470 703520 40582 704960 0 FreeSans 448 90 0 0 io_in[23]
port 44 nsew signal input
flabel metal3 s -960 684164 480 684404 0 FreeSans 960 0 0 0 io_in[24]
port 45 nsew signal input
flabel metal3 s -960 631940 480 632180 0 FreeSans 960 0 0 0 io_in[25]
port 46 nsew signal input
flabel metal3 s -960 579852 480 580092 0 FreeSans 960 0 0 0 io_in[26]
port 47 nsew signal input
flabel metal3 s -960 527764 480 528004 0 FreeSans 960 0 0 0 io_in[27]
port 48 nsew signal input
flabel metal3 s -960 475540 480 475780 0 FreeSans 960 0 0 0 io_in[28]
port 49 nsew signal input
flabel metal3 s -960 423452 480 423692 0 FreeSans 960 0 0 0 io_in[29]
port 50 nsew signal input
flabel metal3 s 583520 86036 584960 86276 0 FreeSans 960 0 0 0 io_in[2]
port 51 nsew signal input
flabel metal3 s -960 371228 480 371468 0 FreeSans 960 0 0 0 io_in[30]
port 52 nsew signal input
flabel metal3 s -960 319140 480 319380 0 FreeSans 960 0 0 0 io_in[31]
port 53 nsew signal input
flabel metal3 s -960 267052 480 267292 0 FreeSans 960 0 0 0 io_in[32]
port 54 nsew signal input
flabel metal3 s -960 214828 480 215068 0 FreeSans 960 0 0 0 io_in[33]
port 55 nsew signal input
flabel metal3 s -960 162740 480 162980 0 FreeSans 960 0 0 0 io_in[34]
port 56 nsew signal input
flabel metal3 s -960 110516 480 110756 0 FreeSans 960 0 0 0 io_in[35]
port 57 nsew signal input
flabel metal3 s -960 71484 480 71724 0 FreeSans 960 0 0 0 io_in[36]
port 58 nsew signal input
flabel metal3 s -960 32316 480 32556 0 FreeSans 960 0 0 0 io_in[37]
port 59 nsew signal input
flabel metal3 s 583520 125884 584960 126124 0 FreeSans 960 0 0 0 io_in[3]
port 60 nsew signal input
flabel metal3 s 583520 165732 584960 165972 0 FreeSans 960 0 0 0 io_in[4]
port 61 nsew signal input
flabel metal3 s 583520 205580 584960 205820 0 FreeSans 960 0 0 0 io_in[5]
port 62 nsew signal input
flabel metal3 s 583520 245428 584960 245668 0 FreeSans 960 0 0 0 io_in[6]
port 63 nsew signal input
flabel metal3 s 583520 298604 584960 298844 0 FreeSans 960 0 0 0 io_in[7]
port 64 nsew signal input
flabel metal3 s 583520 351780 584960 352020 0 FreeSans 960 0 0 0 io_in[8]
port 65 nsew signal input
flabel metal3 s 583520 404820 584960 405060 0 FreeSans 960 0 0 0 io_in[9]
port 66 nsew signal input
flabel metal3 s 583520 32996 584960 33236 0 FreeSans 960 0 0 0 io_oeb[0]
port 67 nsew signal tristate
flabel metal3 s 583520 484516 584960 484756 0 FreeSans 960 0 0 0 io_oeb[10]
port 68 nsew signal tristate
flabel metal3 s 583520 537692 584960 537932 0 FreeSans 960 0 0 0 io_oeb[11]
port 69 nsew signal tristate
flabel metal3 s 583520 590868 584960 591108 0 FreeSans 960 0 0 0 io_oeb[12]
port 70 nsew signal tristate
flabel metal3 s 583520 643908 584960 644148 0 FreeSans 960 0 0 0 io_oeb[13]
port 71 nsew signal tristate
flabel metal3 s 583520 697084 584960 697324 0 FreeSans 960 0 0 0 io_oeb[14]
port 72 nsew signal tristate
flabel metal2 s 527150 703520 527262 704960 0 FreeSans 448 90 0 0 io_oeb[15]
port 73 nsew signal tristate
flabel metal2 s 462290 703520 462402 704960 0 FreeSans 448 90 0 0 io_oeb[16]
port 74 nsew signal tristate
flabel metal2 s 397430 703520 397542 704960 0 FreeSans 448 90 0 0 io_oeb[17]
port 75 nsew signal tristate
flabel metal2 s 332478 703520 332590 704960 0 FreeSans 448 90 0 0 io_oeb[18]
port 76 nsew signal tristate
flabel metal2 s 267618 703520 267730 704960 0 FreeSans 448 90 0 0 io_oeb[19]
port 77 nsew signal tristate
flabel metal3 s 583520 72844 584960 73084 0 FreeSans 960 0 0 0 io_oeb[1]
port 78 nsew signal tristate
flabel metal2 s 202758 703520 202870 704960 0 FreeSans 448 90 0 0 io_oeb[20]
port 79 nsew signal tristate
flabel metal2 s 137806 703520 137918 704960 0 FreeSans 448 90 0 0 io_oeb[21]
port 80 nsew signal tristate
flabel metal2 s 72946 703520 73058 704960 0 FreeSans 448 90 0 0 io_oeb[22]
port 81 nsew signal tristate
flabel metal2 s 8086 703520 8198 704960 0 FreeSans 448 90 0 0 io_oeb[23]
port 82 nsew signal tristate
flabel metal3 s -960 658052 480 658292 0 FreeSans 960 0 0 0 io_oeb[24]
port 83 nsew signal tristate
flabel metal3 s -960 605964 480 606204 0 FreeSans 960 0 0 0 io_oeb[25]
port 84 nsew signal tristate
flabel metal3 s -960 553740 480 553980 0 FreeSans 960 0 0 0 io_oeb[26]
port 85 nsew signal tristate
flabel metal3 s -960 501652 480 501892 0 FreeSans 960 0 0 0 io_oeb[27]
port 86 nsew signal tristate
flabel metal3 s -960 449428 480 449668 0 FreeSans 960 0 0 0 io_oeb[28]
port 87 nsew signal tristate
flabel metal3 s -960 397340 480 397580 0 FreeSans 960 0 0 0 io_oeb[29]
port 88 nsew signal tristate
flabel metal3 s 583520 112692 584960 112932 0 FreeSans 960 0 0 0 io_oeb[2]
port 89 nsew signal tristate
flabel metal3 s -960 345252 480 345492 0 FreeSans 960 0 0 0 io_oeb[30]
port 90 nsew signal tristate
flabel metal3 s -960 293028 480 293268 0 FreeSans 960 0 0 0 io_oeb[31]
port 91 nsew signal tristate
flabel metal3 s -960 240940 480 241180 0 FreeSans 960 0 0 0 io_oeb[32]
port 92 nsew signal tristate
flabel metal3 s -960 188716 480 188956 0 FreeSans 960 0 0 0 io_oeb[33]
port 93 nsew signal tristate
flabel metal3 s -960 136628 480 136868 0 FreeSans 960 0 0 0 io_oeb[34]
port 94 nsew signal tristate
flabel metal3 s -960 84540 480 84780 0 FreeSans 960 0 0 0 io_oeb[35]
port 95 nsew signal tristate
flabel metal3 s -960 45372 480 45612 0 FreeSans 960 0 0 0 io_oeb[36]
port 96 nsew signal tristate
flabel metal3 s -960 6340 480 6580 0 FreeSans 960 0 0 0 io_oeb[37]
port 97 nsew signal tristate
flabel metal3 s 583520 152540 584960 152780 0 FreeSans 960 0 0 0 io_oeb[3]
port 98 nsew signal tristate
flabel metal3 s 583520 192388 584960 192628 0 FreeSans 960 0 0 0 io_oeb[4]
port 99 nsew signal tristate
flabel metal3 s 583520 232236 584960 232476 0 FreeSans 960 0 0 0 io_oeb[5]
port 100 nsew signal tristate
flabel metal3 s 583520 272084 584960 272324 0 FreeSans 960 0 0 0 io_oeb[6]
port 101 nsew signal tristate
flabel metal3 s 583520 325124 584960 325364 0 FreeSans 960 0 0 0 io_oeb[7]
port 102 nsew signal tristate
flabel metal3 s 583520 378300 584960 378540 0 FreeSans 960 0 0 0 io_oeb[8]
port 103 nsew signal tristate
flabel metal3 s 583520 431476 584960 431716 0 FreeSans 960 0 0 0 io_oeb[9]
port 104 nsew signal tristate
flabel metal3 s 583520 19668 584960 19908 0 FreeSans 960 0 0 0 io_out[0]
port 105 nsew signal tristate
flabel metal3 s 583520 471324 584960 471564 0 FreeSans 960 0 0 0 io_out[10]
port 106 nsew signal tristate
flabel metal3 s 583520 524364 584960 524604 0 FreeSans 960 0 0 0 io_out[11]
port 107 nsew signal tristate
flabel metal3 s 583520 577540 584960 577780 0 FreeSans 960 0 0 0 io_out[12]
port 108 nsew signal tristate
flabel metal3 s 583520 630716 584960 630956 0 FreeSans 960 0 0 0 io_out[13]
port 109 nsew signal tristate
flabel metal3 s 583520 683756 584960 683996 0 FreeSans 960 0 0 0 io_out[14]
port 110 nsew signal tristate
flabel metal2 s 543434 703520 543546 704960 0 FreeSans 448 90 0 0 io_out[15]
port 111 nsew signal tristate
flabel metal2 s 478482 703520 478594 704960 0 FreeSans 448 90 0 0 io_out[16]
port 112 nsew signal tristate
flabel metal2 s 413622 703520 413734 704960 0 FreeSans 448 90 0 0 io_out[17]
port 113 nsew signal tristate
flabel metal2 s 348762 703520 348874 704960 0 FreeSans 448 90 0 0 io_out[18]
port 114 nsew signal tristate
flabel metal2 s 283810 703520 283922 704960 0 FreeSans 448 90 0 0 io_out[19]
port 115 nsew signal tristate
flabel metal3 s 583520 59516 584960 59756 0 FreeSans 960 0 0 0 io_out[1]
port 116 nsew signal tristate
flabel metal2 s 218950 703520 219062 704960 0 FreeSans 448 90 0 0 io_out[20]
port 117 nsew signal tristate
flabel metal2 s 154090 703520 154202 704960 0 FreeSans 448 90 0 0 io_out[21]
port 118 nsew signal tristate
flabel metal2 s 89138 703520 89250 704960 0 FreeSans 448 90 0 0 io_out[22]
port 119 nsew signal tristate
flabel metal2 s 24278 703520 24390 704960 0 FreeSans 448 90 0 0 io_out[23]
port 120 nsew signal tristate
flabel metal3 s -960 671108 480 671348 0 FreeSans 960 0 0 0 io_out[24]
port 121 nsew signal tristate
flabel metal3 s -960 619020 480 619260 0 FreeSans 960 0 0 0 io_out[25]
port 122 nsew signal tristate
flabel metal3 s -960 566796 480 567036 0 FreeSans 960 0 0 0 io_out[26]
port 123 nsew signal tristate
flabel metal3 s -960 514708 480 514948 0 FreeSans 960 0 0 0 io_out[27]
port 124 nsew signal tristate
flabel metal3 s -960 462484 480 462724 0 FreeSans 960 0 0 0 io_out[28]
port 125 nsew signal tristate
flabel metal3 s -960 410396 480 410636 0 FreeSans 960 0 0 0 io_out[29]
port 126 nsew signal tristate
flabel metal3 s 583520 99364 584960 99604 0 FreeSans 960 0 0 0 io_out[2]
port 127 nsew signal tristate
flabel metal3 s -960 358308 480 358548 0 FreeSans 960 0 0 0 io_out[30]
port 128 nsew signal tristate
flabel metal3 s -960 306084 480 306324 0 FreeSans 960 0 0 0 io_out[31]
port 129 nsew signal tristate
flabel metal3 s -960 253996 480 254236 0 FreeSans 960 0 0 0 io_out[32]
port 130 nsew signal tristate
flabel metal3 s -960 201772 480 202012 0 FreeSans 960 0 0 0 io_out[33]
port 131 nsew signal tristate
flabel metal3 s -960 149684 480 149924 0 FreeSans 960 0 0 0 io_out[34]
port 132 nsew signal tristate
flabel metal3 s -960 97460 480 97700 0 FreeSans 960 0 0 0 io_out[35]
port 133 nsew signal tristate
flabel metal3 s -960 58428 480 58668 0 FreeSans 960 0 0 0 io_out[36]
port 134 nsew signal tristate
flabel metal3 s -960 19260 480 19500 0 FreeSans 960 0 0 0 io_out[37]
port 135 nsew signal tristate
flabel metal3 s 583520 139212 584960 139452 0 FreeSans 960 0 0 0 io_out[3]
port 136 nsew signal tristate
flabel metal3 s 583520 179060 584960 179300 0 FreeSans 960 0 0 0 io_out[4]
port 137 nsew signal tristate
flabel metal3 s 583520 218908 584960 219148 0 FreeSans 960 0 0 0 io_out[5]
port 138 nsew signal tristate
flabel metal3 s 583520 258756 584960 258996 0 FreeSans 960 0 0 0 io_out[6]
port 139 nsew signal tristate
flabel metal3 s 583520 311932 584960 312172 0 FreeSans 960 0 0 0 io_out[7]
port 140 nsew signal tristate
flabel metal3 s 583520 364972 584960 365212 0 FreeSans 960 0 0 0 io_out[8]
port 141 nsew signal tristate
flabel metal3 s 583520 418148 584960 418388 0 FreeSans 960 0 0 0 io_out[9]
port 142 nsew signal tristate
flabel metal2 s 125846 -960 125958 480 0 FreeSans 448 90 0 0 la_data_in[0]
port 143 nsew signal input
flabel metal2 s 480506 -960 480618 480 0 FreeSans 448 90 0 0 la_data_in[100]
port 144 nsew signal input
flabel metal2 s 484002 -960 484114 480 0 FreeSans 448 90 0 0 la_data_in[101]
port 145 nsew signal input
flabel metal2 s 487590 -960 487702 480 0 FreeSans 448 90 0 0 la_data_in[102]
port 146 nsew signal input
flabel metal2 s 491086 -960 491198 480 0 FreeSans 448 90 0 0 la_data_in[103]
port 147 nsew signal input
flabel metal2 s 494674 -960 494786 480 0 FreeSans 448 90 0 0 la_data_in[104]
port 148 nsew signal input
flabel metal2 s 498170 -960 498282 480 0 FreeSans 448 90 0 0 la_data_in[105]
port 149 nsew signal input
flabel metal2 s 501758 -960 501870 480 0 FreeSans 448 90 0 0 la_data_in[106]
port 150 nsew signal input
flabel metal2 s 505346 -960 505458 480 0 FreeSans 448 90 0 0 la_data_in[107]
port 151 nsew signal input
flabel metal2 s 508842 -960 508954 480 0 FreeSans 448 90 0 0 la_data_in[108]
port 152 nsew signal input
flabel metal2 s 512430 -960 512542 480 0 FreeSans 448 90 0 0 la_data_in[109]
port 153 nsew signal input
flabel metal2 s 161266 -960 161378 480 0 FreeSans 448 90 0 0 la_data_in[10]
port 154 nsew signal input
flabel metal2 s 515926 -960 516038 480 0 FreeSans 448 90 0 0 la_data_in[110]
port 155 nsew signal input
flabel metal2 s 519514 -960 519626 480 0 FreeSans 448 90 0 0 la_data_in[111]
port 156 nsew signal input
flabel metal2 s 523010 -960 523122 480 0 FreeSans 448 90 0 0 la_data_in[112]
port 157 nsew signal input
flabel metal2 s 526598 -960 526710 480 0 FreeSans 448 90 0 0 la_data_in[113]
port 158 nsew signal input
flabel metal2 s 530094 -960 530206 480 0 FreeSans 448 90 0 0 la_data_in[114]
port 159 nsew signal input
flabel metal2 s 533682 -960 533794 480 0 FreeSans 448 90 0 0 la_data_in[115]
port 160 nsew signal input
flabel metal2 s 537178 -960 537290 480 0 FreeSans 448 90 0 0 la_data_in[116]
port 161 nsew signal input
flabel metal2 s 540766 -960 540878 480 0 FreeSans 448 90 0 0 la_data_in[117]
port 162 nsew signal input
flabel metal2 s 544354 -960 544466 480 0 FreeSans 448 90 0 0 la_data_in[118]
port 163 nsew signal input
flabel metal2 s 547850 -960 547962 480 0 FreeSans 448 90 0 0 la_data_in[119]
port 164 nsew signal input
flabel metal2 s 164854 -960 164966 480 0 FreeSans 448 90 0 0 la_data_in[11]
port 165 nsew signal input
flabel metal2 s 551438 -960 551550 480 0 FreeSans 448 90 0 0 la_data_in[120]
port 166 nsew signal input
flabel metal2 s 554934 -960 555046 480 0 FreeSans 448 90 0 0 la_data_in[121]
port 167 nsew signal input
flabel metal2 s 558522 -960 558634 480 0 FreeSans 448 90 0 0 la_data_in[122]
port 168 nsew signal input
flabel metal2 s 562018 -960 562130 480 0 FreeSans 448 90 0 0 la_data_in[123]
port 169 nsew signal input
flabel metal2 s 565606 -960 565718 480 0 FreeSans 448 90 0 0 la_data_in[124]
port 170 nsew signal input
flabel metal2 s 569102 -960 569214 480 0 FreeSans 448 90 0 0 la_data_in[125]
port 171 nsew signal input
flabel metal2 s 572690 -960 572802 480 0 FreeSans 448 90 0 0 la_data_in[126]
port 172 nsew signal input
flabel metal2 s 576278 -960 576390 480 0 FreeSans 448 90 0 0 la_data_in[127]
port 173 nsew signal input
flabel metal2 s 168350 -960 168462 480 0 FreeSans 448 90 0 0 la_data_in[12]
port 174 nsew signal input
flabel metal2 s 171938 -960 172050 480 0 FreeSans 448 90 0 0 la_data_in[13]
port 175 nsew signal input
flabel metal2 s 175434 -960 175546 480 0 FreeSans 448 90 0 0 la_data_in[14]
port 176 nsew signal input
flabel metal2 s 179022 -960 179134 480 0 FreeSans 448 90 0 0 la_data_in[15]
port 177 nsew signal input
flabel metal2 s 182518 -960 182630 480 0 FreeSans 448 90 0 0 la_data_in[16]
port 178 nsew signal input
flabel metal2 s 186106 -960 186218 480 0 FreeSans 448 90 0 0 la_data_in[17]
port 179 nsew signal input
flabel metal2 s 189694 -960 189806 480 0 FreeSans 448 90 0 0 la_data_in[18]
port 180 nsew signal input
flabel metal2 s 193190 -960 193302 480 0 FreeSans 448 90 0 0 la_data_in[19]
port 181 nsew signal input
flabel metal2 s 129342 -960 129454 480 0 FreeSans 448 90 0 0 la_data_in[1]
port 182 nsew signal input
flabel metal2 s 196778 -960 196890 480 0 FreeSans 448 90 0 0 la_data_in[20]
port 183 nsew signal input
flabel metal2 s 200274 -960 200386 480 0 FreeSans 448 90 0 0 la_data_in[21]
port 184 nsew signal input
flabel metal2 s 203862 -960 203974 480 0 FreeSans 448 90 0 0 la_data_in[22]
port 185 nsew signal input
flabel metal2 s 207358 -960 207470 480 0 FreeSans 448 90 0 0 la_data_in[23]
port 186 nsew signal input
flabel metal2 s 210946 -960 211058 480 0 FreeSans 448 90 0 0 la_data_in[24]
port 187 nsew signal input
flabel metal2 s 214442 -960 214554 480 0 FreeSans 448 90 0 0 la_data_in[25]
port 188 nsew signal input
flabel metal2 s 218030 -960 218142 480 0 FreeSans 448 90 0 0 la_data_in[26]
port 189 nsew signal input
flabel metal2 s 221526 -960 221638 480 0 FreeSans 448 90 0 0 la_data_in[27]
port 190 nsew signal input
flabel metal2 s 225114 -960 225226 480 0 FreeSans 448 90 0 0 la_data_in[28]
port 191 nsew signal input
flabel metal2 s 228702 -960 228814 480 0 FreeSans 448 90 0 0 la_data_in[29]
port 192 nsew signal input
flabel metal2 s 132930 -960 133042 480 0 FreeSans 448 90 0 0 la_data_in[2]
port 193 nsew signal input
flabel metal2 s 232198 -960 232310 480 0 FreeSans 448 90 0 0 la_data_in[30]
port 194 nsew signal input
flabel metal2 s 235786 -960 235898 480 0 FreeSans 448 90 0 0 la_data_in[31]
port 195 nsew signal input
flabel metal2 s 239282 -960 239394 480 0 FreeSans 448 90 0 0 la_data_in[32]
port 196 nsew signal input
flabel metal2 s 242870 -960 242982 480 0 FreeSans 448 90 0 0 la_data_in[33]
port 197 nsew signal input
flabel metal2 s 246366 -960 246478 480 0 FreeSans 448 90 0 0 la_data_in[34]
port 198 nsew signal input
flabel metal2 s 249954 -960 250066 480 0 FreeSans 448 90 0 0 la_data_in[35]
port 199 nsew signal input
flabel metal2 s 253450 -960 253562 480 0 FreeSans 448 90 0 0 la_data_in[36]
port 200 nsew signal input
flabel metal2 s 257038 -960 257150 480 0 FreeSans 448 90 0 0 la_data_in[37]
port 201 nsew signal input
flabel metal2 s 260626 -960 260738 480 0 FreeSans 448 90 0 0 la_data_in[38]
port 202 nsew signal input
flabel metal2 s 264122 -960 264234 480 0 FreeSans 448 90 0 0 la_data_in[39]
port 203 nsew signal input
flabel metal2 s 136426 -960 136538 480 0 FreeSans 448 90 0 0 la_data_in[3]
port 204 nsew signal input
flabel metal2 s 267710 -960 267822 480 0 FreeSans 448 90 0 0 la_data_in[40]
port 205 nsew signal input
flabel metal2 s 271206 -960 271318 480 0 FreeSans 448 90 0 0 la_data_in[41]
port 206 nsew signal input
flabel metal2 s 274794 -960 274906 480 0 FreeSans 448 90 0 0 la_data_in[42]
port 207 nsew signal input
flabel metal2 s 278290 -960 278402 480 0 FreeSans 448 90 0 0 la_data_in[43]
port 208 nsew signal input
flabel metal2 s 281878 -960 281990 480 0 FreeSans 448 90 0 0 la_data_in[44]
port 209 nsew signal input
flabel metal2 s 285374 -960 285486 480 0 FreeSans 448 90 0 0 la_data_in[45]
port 210 nsew signal input
flabel metal2 s 288962 -960 289074 480 0 FreeSans 448 90 0 0 la_data_in[46]
port 211 nsew signal input
flabel metal2 s 292550 -960 292662 480 0 FreeSans 448 90 0 0 la_data_in[47]
port 212 nsew signal input
flabel metal2 s 296046 -960 296158 480 0 FreeSans 448 90 0 0 la_data_in[48]
port 213 nsew signal input
flabel metal2 s 299634 -960 299746 480 0 FreeSans 448 90 0 0 la_data_in[49]
port 214 nsew signal input
flabel metal2 s 140014 -960 140126 480 0 FreeSans 448 90 0 0 la_data_in[4]
port 215 nsew signal input
flabel metal2 s 303130 -960 303242 480 0 FreeSans 448 90 0 0 la_data_in[50]
port 216 nsew signal input
flabel metal2 s 306718 -960 306830 480 0 FreeSans 448 90 0 0 la_data_in[51]
port 217 nsew signal input
flabel metal2 s 310214 -960 310326 480 0 FreeSans 448 90 0 0 la_data_in[52]
port 218 nsew signal input
flabel metal2 s 313802 -960 313914 480 0 FreeSans 448 90 0 0 la_data_in[53]
port 219 nsew signal input
flabel metal2 s 317298 -960 317410 480 0 FreeSans 448 90 0 0 la_data_in[54]
port 220 nsew signal input
flabel metal2 s 320886 -960 320998 480 0 FreeSans 448 90 0 0 la_data_in[55]
port 221 nsew signal input
flabel metal2 s 324382 -960 324494 480 0 FreeSans 448 90 0 0 la_data_in[56]
port 222 nsew signal input
flabel metal2 s 327970 -960 328082 480 0 FreeSans 448 90 0 0 la_data_in[57]
port 223 nsew signal input
flabel metal2 s 331558 -960 331670 480 0 FreeSans 448 90 0 0 la_data_in[58]
port 224 nsew signal input
flabel metal2 s 335054 -960 335166 480 0 FreeSans 448 90 0 0 la_data_in[59]
port 225 nsew signal input
flabel metal2 s 143510 -960 143622 480 0 FreeSans 448 90 0 0 la_data_in[5]
port 226 nsew signal input
flabel metal2 s 338642 -960 338754 480 0 FreeSans 448 90 0 0 la_data_in[60]
port 227 nsew signal input
flabel metal2 s 342138 -960 342250 480 0 FreeSans 448 90 0 0 la_data_in[61]
port 228 nsew signal input
flabel metal2 s 345726 -960 345838 480 0 FreeSans 448 90 0 0 la_data_in[62]
port 229 nsew signal input
flabel metal2 s 349222 -960 349334 480 0 FreeSans 448 90 0 0 la_data_in[63]
port 230 nsew signal input
flabel metal2 s 352810 -960 352922 480 0 FreeSans 448 90 0 0 la_data_in[64]
port 231 nsew signal input
flabel metal2 s 356306 -960 356418 480 0 FreeSans 448 90 0 0 la_data_in[65]
port 232 nsew signal input
flabel metal2 s 359894 -960 360006 480 0 FreeSans 448 90 0 0 la_data_in[66]
port 233 nsew signal input
flabel metal2 s 363482 -960 363594 480 0 FreeSans 448 90 0 0 la_data_in[67]
port 234 nsew signal input
flabel metal2 s 366978 -960 367090 480 0 FreeSans 448 90 0 0 la_data_in[68]
port 235 nsew signal input
flabel metal2 s 370566 -960 370678 480 0 FreeSans 448 90 0 0 la_data_in[69]
port 236 nsew signal input
flabel metal2 s 147098 -960 147210 480 0 FreeSans 448 90 0 0 la_data_in[6]
port 237 nsew signal input
flabel metal2 s 374062 -960 374174 480 0 FreeSans 448 90 0 0 la_data_in[70]
port 238 nsew signal input
flabel metal2 s 377650 -960 377762 480 0 FreeSans 448 90 0 0 la_data_in[71]
port 239 nsew signal input
flabel metal2 s 381146 -960 381258 480 0 FreeSans 448 90 0 0 la_data_in[72]
port 240 nsew signal input
flabel metal2 s 384734 -960 384846 480 0 FreeSans 448 90 0 0 la_data_in[73]
port 241 nsew signal input
flabel metal2 s 388230 -960 388342 480 0 FreeSans 448 90 0 0 la_data_in[74]
port 242 nsew signal input
flabel metal2 s 391818 -960 391930 480 0 FreeSans 448 90 0 0 la_data_in[75]
port 243 nsew signal input
flabel metal2 s 395314 -960 395426 480 0 FreeSans 448 90 0 0 la_data_in[76]
port 244 nsew signal input
flabel metal2 s 398902 -960 399014 480 0 FreeSans 448 90 0 0 la_data_in[77]
port 245 nsew signal input
flabel metal2 s 402490 -960 402602 480 0 FreeSans 448 90 0 0 la_data_in[78]
port 246 nsew signal input
flabel metal2 s 405986 -960 406098 480 0 FreeSans 448 90 0 0 la_data_in[79]
port 247 nsew signal input
flabel metal2 s 150594 -960 150706 480 0 FreeSans 448 90 0 0 la_data_in[7]
port 248 nsew signal input
flabel metal2 s 409574 -960 409686 480 0 FreeSans 448 90 0 0 la_data_in[80]
port 249 nsew signal input
flabel metal2 s 413070 -960 413182 480 0 FreeSans 448 90 0 0 la_data_in[81]
port 250 nsew signal input
flabel metal2 s 416658 -960 416770 480 0 FreeSans 448 90 0 0 la_data_in[82]
port 251 nsew signal input
flabel metal2 s 420154 -960 420266 480 0 FreeSans 448 90 0 0 la_data_in[83]
port 252 nsew signal input
flabel metal2 s 423742 -960 423854 480 0 FreeSans 448 90 0 0 la_data_in[84]
port 253 nsew signal input
flabel metal2 s 427238 -960 427350 480 0 FreeSans 448 90 0 0 la_data_in[85]
port 254 nsew signal input
flabel metal2 s 430826 -960 430938 480 0 FreeSans 448 90 0 0 la_data_in[86]
port 255 nsew signal input
flabel metal2 s 434414 -960 434526 480 0 FreeSans 448 90 0 0 la_data_in[87]
port 256 nsew signal input
flabel metal2 s 437910 -960 438022 480 0 FreeSans 448 90 0 0 la_data_in[88]
port 257 nsew signal input
flabel metal2 s 441498 -960 441610 480 0 FreeSans 448 90 0 0 la_data_in[89]
port 258 nsew signal input
flabel metal2 s 154182 -960 154294 480 0 FreeSans 448 90 0 0 la_data_in[8]
port 259 nsew signal input
flabel metal2 s 444994 -960 445106 480 0 FreeSans 448 90 0 0 la_data_in[90]
port 260 nsew signal input
flabel metal2 s 448582 -960 448694 480 0 FreeSans 448 90 0 0 la_data_in[91]
port 261 nsew signal input
flabel metal2 s 452078 -960 452190 480 0 FreeSans 448 90 0 0 la_data_in[92]
port 262 nsew signal input
flabel metal2 s 455666 -960 455778 480 0 FreeSans 448 90 0 0 la_data_in[93]
port 263 nsew signal input
flabel metal2 s 459162 -960 459274 480 0 FreeSans 448 90 0 0 la_data_in[94]
port 264 nsew signal input
flabel metal2 s 462750 -960 462862 480 0 FreeSans 448 90 0 0 la_data_in[95]
port 265 nsew signal input
flabel metal2 s 466246 -960 466358 480 0 FreeSans 448 90 0 0 la_data_in[96]
port 266 nsew signal input
flabel metal2 s 469834 -960 469946 480 0 FreeSans 448 90 0 0 la_data_in[97]
port 267 nsew signal input
flabel metal2 s 473422 -960 473534 480 0 FreeSans 448 90 0 0 la_data_in[98]
port 268 nsew signal input
flabel metal2 s 476918 -960 477030 480 0 FreeSans 448 90 0 0 la_data_in[99]
port 269 nsew signal input
flabel metal2 s 157770 -960 157882 480 0 FreeSans 448 90 0 0 la_data_in[9]
port 270 nsew signal input
flabel metal2 s 126950 -960 127062 480 0 FreeSans 448 90 0 0 la_data_out[0]
port 271 nsew signal tristate
flabel metal2 s 481702 -960 481814 480 0 FreeSans 448 90 0 0 la_data_out[100]
port 272 nsew signal tristate
flabel metal2 s 485198 -960 485310 480 0 FreeSans 448 90 0 0 la_data_out[101]
port 273 nsew signal tristate
flabel metal2 s 488786 -960 488898 480 0 FreeSans 448 90 0 0 la_data_out[102]
port 274 nsew signal tristate
flabel metal2 s 492282 -960 492394 480 0 FreeSans 448 90 0 0 la_data_out[103]
port 275 nsew signal tristate
flabel metal2 s 495870 -960 495982 480 0 FreeSans 448 90 0 0 la_data_out[104]
port 276 nsew signal tristate
flabel metal2 s 499366 -960 499478 480 0 FreeSans 448 90 0 0 la_data_out[105]
port 277 nsew signal tristate
flabel metal2 s 502954 -960 503066 480 0 FreeSans 448 90 0 0 la_data_out[106]
port 278 nsew signal tristate
flabel metal2 s 506450 -960 506562 480 0 FreeSans 448 90 0 0 la_data_out[107]
port 279 nsew signal tristate
flabel metal2 s 510038 -960 510150 480 0 FreeSans 448 90 0 0 la_data_out[108]
port 280 nsew signal tristate
flabel metal2 s 513534 -960 513646 480 0 FreeSans 448 90 0 0 la_data_out[109]
port 281 nsew signal tristate
flabel metal2 s 162462 -960 162574 480 0 FreeSans 448 90 0 0 la_data_out[10]
port 282 nsew signal tristate
flabel metal2 s 517122 -960 517234 480 0 FreeSans 448 90 0 0 la_data_out[110]
port 283 nsew signal tristate
flabel metal2 s 520710 -960 520822 480 0 FreeSans 448 90 0 0 la_data_out[111]
port 284 nsew signal tristate
flabel metal2 s 524206 -960 524318 480 0 FreeSans 448 90 0 0 la_data_out[112]
port 285 nsew signal tristate
flabel metal2 s 527794 -960 527906 480 0 FreeSans 448 90 0 0 la_data_out[113]
port 286 nsew signal tristate
flabel metal2 s 531290 -960 531402 480 0 FreeSans 448 90 0 0 la_data_out[114]
port 287 nsew signal tristate
flabel metal2 s 534878 -960 534990 480 0 FreeSans 448 90 0 0 la_data_out[115]
port 288 nsew signal tristate
flabel metal2 s 538374 -960 538486 480 0 FreeSans 448 90 0 0 la_data_out[116]
port 289 nsew signal tristate
flabel metal2 s 541962 -960 542074 480 0 FreeSans 448 90 0 0 la_data_out[117]
port 290 nsew signal tristate
flabel metal2 s 545458 -960 545570 480 0 FreeSans 448 90 0 0 la_data_out[118]
port 291 nsew signal tristate
flabel metal2 s 549046 -960 549158 480 0 FreeSans 448 90 0 0 la_data_out[119]
port 292 nsew signal tristate
flabel metal2 s 166050 -960 166162 480 0 FreeSans 448 90 0 0 la_data_out[11]
port 293 nsew signal tristate
flabel metal2 s 552634 -960 552746 480 0 FreeSans 448 90 0 0 la_data_out[120]
port 294 nsew signal tristate
flabel metal2 s 556130 -960 556242 480 0 FreeSans 448 90 0 0 la_data_out[121]
port 295 nsew signal tristate
flabel metal2 s 559718 -960 559830 480 0 FreeSans 448 90 0 0 la_data_out[122]
port 296 nsew signal tristate
flabel metal2 s 563214 -960 563326 480 0 FreeSans 448 90 0 0 la_data_out[123]
port 297 nsew signal tristate
flabel metal2 s 566802 -960 566914 480 0 FreeSans 448 90 0 0 la_data_out[124]
port 298 nsew signal tristate
flabel metal2 s 570298 -960 570410 480 0 FreeSans 448 90 0 0 la_data_out[125]
port 299 nsew signal tristate
flabel metal2 s 573886 -960 573998 480 0 FreeSans 448 90 0 0 la_data_out[126]
port 300 nsew signal tristate
flabel metal2 s 577382 -960 577494 480 0 FreeSans 448 90 0 0 la_data_out[127]
port 301 nsew signal tristate
flabel metal2 s 169546 -960 169658 480 0 FreeSans 448 90 0 0 la_data_out[12]
port 302 nsew signal tristate
flabel metal2 s 173134 -960 173246 480 0 FreeSans 448 90 0 0 la_data_out[13]
port 303 nsew signal tristate
flabel metal2 s 176630 -960 176742 480 0 FreeSans 448 90 0 0 la_data_out[14]
port 304 nsew signal tristate
flabel metal2 s 180218 -960 180330 480 0 FreeSans 448 90 0 0 la_data_out[15]
port 305 nsew signal tristate
flabel metal2 s 183714 -960 183826 480 0 FreeSans 448 90 0 0 la_data_out[16]
port 306 nsew signal tristate
flabel metal2 s 187302 -960 187414 480 0 FreeSans 448 90 0 0 la_data_out[17]
port 307 nsew signal tristate
flabel metal2 s 190798 -960 190910 480 0 FreeSans 448 90 0 0 la_data_out[18]
port 308 nsew signal tristate
flabel metal2 s 194386 -960 194498 480 0 FreeSans 448 90 0 0 la_data_out[19]
port 309 nsew signal tristate
flabel metal2 s 130538 -960 130650 480 0 FreeSans 448 90 0 0 la_data_out[1]
port 310 nsew signal tristate
flabel metal2 s 197882 -960 197994 480 0 FreeSans 448 90 0 0 la_data_out[20]
port 311 nsew signal tristate
flabel metal2 s 201470 -960 201582 480 0 FreeSans 448 90 0 0 la_data_out[21]
port 312 nsew signal tristate
flabel metal2 s 205058 -960 205170 480 0 FreeSans 448 90 0 0 la_data_out[22]
port 313 nsew signal tristate
flabel metal2 s 208554 -960 208666 480 0 FreeSans 448 90 0 0 la_data_out[23]
port 314 nsew signal tristate
flabel metal2 s 212142 -960 212254 480 0 FreeSans 448 90 0 0 la_data_out[24]
port 315 nsew signal tristate
flabel metal2 s 215638 -960 215750 480 0 FreeSans 448 90 0 0 la_data_out[25]
port 316 nsew signal tristate
flabel metal2 s 219226 -960 219338 480 0 FreeSans 448 90 0 0 la_data_out[26]
port 317 nsew signal tristate
flabel metal2 s 222722 -960 222834 480 0 FreeSans 448 90 0 0 la_data_out[27]
port 318 nsew signal tristate
flabel metal2 s 226310 -960 226422 480 0 FreeSans 448 90 0 0 la_data_out[28]
port 319 nsew signal tristate
flabel metal2 s 229806 -960 229918 480 0 FreeSans 448 90 0 0 la_data_out[29]
port 320 nsew signal tristate
flabel metal2 s 134126 -960 134238 480 0 FreeSans 448 90 0 0 la_data_out[2]
port 321 nsew signal tristate
flabel metal2 s 233394 -960 233506 480 0 FreeSans 448 90 0 0 la_data_out[30]
port 322 nsew signal tristate
flabel metal2 s 236982 -960 237094 480 0 FreeSans 448 90 0 0 la_data_out[31]
port 323 nsew signal tristate
flabel metal2 s 240478 -960 240590 480 0 FreeSans 448 90 0 0 la_data_out[32]
port 324 nsew signal tristate
flabel metal2 s 244066 -960 244178 480 0 FreeSans 448 90 0 0 la_data_out[33]
port 325 nsew signal tristate
flabel metal2 s 247562 -960 247674 480 0 FreeSans 448 90 0 0 la_data_out[34]
port 326 nsew signal tristate
flabel metal2 s 251150 -960 251262 480 0 FreeSans 448 90 0 0 la_data_out[35]
port 327 nsew signal tristate
flabel metal2 s 254646 -960 254758 480 0 FreeSans 448 90 0 0 la_data_out[36]
port 328 nsew signal tristate
flabel metal2 s 258234 -960 258346 480 0 FreeSans 448 90 0 0 la_data_out[37]
port 329 nsew signal tristate
flabel metal2 s 261730 -960 261842 480 0 FreeSans 448 90 0 0 la_data_out[38]
port 330 nsew signal tristate
flabel metal2 s 265318 -960 265430 480 0 FreeSans 448 90 0 0 la_data_out[39]
port 331 nsew signal tristate
flabel metal2 s 137622 -960 137734 480 0 FreeSans 448 90 0 0 la_data_out[3]
port 332 nsew signal tristate
flabel metal2 s 268814 -960 268926 480 0 FreeSans 448 90 0 0 la_data_out[40]
port 333 nsew signal tristate
flabel metal2 s 272402 -960 272514 480 0 FreeSans 448 90 0 0 la_data_out[41]
port 334 nsew signal tristate
flabel metal2 s 275990 -960 276102 480 0 FreeSans 448 90 0 0 la_data_out[42]
port 335 nsew signal tristate
flabel metal2 s 279486 -960 279598 480 0 FreeSans 448 90 0 0 la_data_out[43]
port 336 nsew signal tristate
flabel metal2 s 283074 -960 283186 480 0 FreeSans 448 90 0 0 la_data_out[44]
port 337 nsew signal tristate
flabel metal2 s 286570 -960 286682 480 0 FreeSans 448 90 0 0 la_data_out[45]
port 338 nsew signal tristate
flabel metal2 s 290158 -960 290270 480 0 FreeSans 448 90 0 0 la_data_out[46]
port 339 nsew signal tristate
flabel metal2 s 293654 -960 293766 480 0 FreeSans 448 90 0 0 la_data_out[47]
port 340 nsew signal tristate
flabel metal2 s 297242 -960 297354 480 0 FreeSans 448 90 0 0 la_data_out[48]
port 341 nsew signal tristate
flabel metal2 s 300738 -960 300850 480 0 FreeSans 448 90 0 0 la_data_out[49]
port 342 nsew signal tristate
flabel metal2 s 141210 -960 141322 480 0 FreeSans 448 90 0 0 la_data_out[4]
port 343 nsew signal tristate
flabel metal2 s 304326 -960 304438 480 0 FreeSans 448 90 0 0 la_data_out[50]
port 344 nsew signal tristate
flabel metal2 s 307914 -960 308026 480 0 FreeSans 448 90 0 0 la_data_out[51]
port 345 nsew signal tristate
flabel metal2 s 311410 -960 311522 480 0 FreeSans 448 90 0 0 la_data_out[52]
port 346 nsew signal tristate
flabel metal2 s 314998 -960 315110 480 0 FreeSans 448 90 0 0 la_data_out[53]
port 347 nsew signal tristate
flabel metal2 s 318494 -960 318606 480 0 FreeSans 448 90 0 0 la_data_out[54]
port 348 nsew signal tristate
flabel metal2 s 322082 -960 322194 480 0 FreeSans 448 90 0 0 la_data_out[55]
port 349 nsew signal tristate
flabel metal2 s 325578 -960 325690 480 0 FreeSans 448 90 0 0 la_data_out[56]
port 350 nsew signal tristate
flabel metal2 s 329166 -960 329278 480 0 FreeSans 448 90 0 0 la_data_out[57]
port 351 nsew signal tristate
flabel metal2 s 332662 -960 332774 480 0 FreeSans 448 90 0 0 la_data_out[58]
port 352 nsew signal tristate
flabel metal2 s 336250 -960 336362 480 0 FreeSans 448 90 0 0 la_data_out[59]
port 353 nsew signal tristate
flabel metal2 s 144706 -960 144818 480 0 FreeSans 448 90 0 0 la_data_out[5]
port 354 nsew signal tristate
flabel metal2 s 339838 -960 339950 480 0 FreeSans 448 90 0 0 la_data_out[60]
port 355 nsew signal tristate
flabel metal2 s 343334 -960 343446 480 0 FreeSans 448 90 0 0 la_data_out[61]
port 356 nsew signal tristate
flabel metal2 s 346922 -960 347034 480 0 FreeSans 448 90 0 0 la_data_out[62]
port 357 nsew signal tristate
flabel metal2 s 350418 -960 350530 480 0 FreeSans 448 90 0 0 la_data_out[63]
port 358 nsew signal tristate
flabel metal2 s 354006 -960 354118 480 0 FreeSans 448 90 0 0 la_data_out[64]
port 359 nsew signal tristate
flabel metal2 s 357502 -960 357614 480 0 FreeSans 448 90 0 0 la_data_out[65]
port 360 nsew signal tristate
flabel metal2 s 361090 -960 361202 480 0 FreeSans 448 90 0 0 la_data_out[66]
port 361 nsew signal tristate
flabel metal2 s 364586 -960 364698 480 0 FreeSans 448 90 0 0 la_data_out[67]
port 362 nsew signal tristate
flabel metal2 s 368174 -960 368286 480 0 FreeSans 448 90 0 0 la_data_out[68]
port 363 nsew signal tristate
flabel metal2 s 371670 -960 371782 480 0 FreeSans 448 90 0 0 la_data_out[69]
port 364 nsew signal tristate
flabel metal2 s 148294 -960 148406 480 0 FreeSans 448 90 0 0 la_data_out[6]
port 365 nsew signal tristate
flabel metal2 s 375258 -960 375370 480 0 FreeSans 448 90 0 0 la_data_out[70]
port 366 nsew signal tristate
flabel metal2 s 378846 -960 378958 480 0 FreeSans 448 90 0 0 la_data_out[71]
port 367 nsew signal tristate
flabel metal2 s 382342 -960 382454 480 0 FreeSans 448 90 0 0 la_data_out[72]
port 368 nsew signal tristate
flabel metal2 s 385930 -960 386042 480 0 FreeSans 448 90 0 0 la_data_out[73]
port 369 nsew signal tristate
flabel metal2 s 389426 -960 389538 480 0 FreeSans 448 90 0 0 la_data_out[74]
port 370 nsew signal tristate
flabel metal2 s 393014 -960 393126 480 0 FreeSans 448 90 0 0 la_data_out[75]
port 371 nsew signal tristate
flabel metal2 s 396510 -960 396622 480 0 FreeSans 448 90 0 0 la_data_out[76]
port 372 nsew signal tristate
flabel metal2 s 400098 -960 400210 480 0 FreeSans 448 90 0 0 la_data_out[77]
port 373 nsew signal tristate
flabel metal2 s 403594 -960 403706 480 0 FreeSans 448 90 0 0 la_data_out[78]
port 374 nsew signal tristate
flabel metal2 s 407182 -960 407294 480 0 FreeSans 448 90 0 0 la_data_out[79]
port 375 nsew signal tristate
flabel metal2 s 151790 -960 151902 480 0 FreeSans 448 90 0 0 la_data_out[7]
port 376 nsew signal tristate
flabel metal2 s 410770 -960 410882 480 0 FreeSans 448 90 0 0 la_data_out[80]
port 377 nsew signal tristate
flabel metal2 s 414266 -960 414378 480 0 FreeSans 448 90 0 0 la_data_out[81]
port 378 nsew signal tristate
flabel metal2 s 417854 -960 417966 480 0 FreeSans 448 90 0 0 la_data_out[82]
port 379 nsew signal tristate
flabel metal2 s 421350 -960 421462 480 0 FreeSans 448 90 0 0 la_data_out[83]
port 380 nsew signal tristate
flabel metal2 s 424938 -960 425050 480 0 FreeSans 448 90 0 0 la_data_out[84]
port 381 nsew signal tristate
flabel metal2 s 428434 -960 428546 480 0 FreeSans 448 90 0 0 la_data_out[85]
port 382 nsew signal tristate
flabel metal2 s 432022 -960 432134 480 0 FreeSans 448 90 0 0 la_data_out[86]
port 383 nsew signal tristate
flabel metal2 s 435518 -960 435630 480 0 FreeSans 448 90 0 0 la_data_out[87]
port 384 nsew signal tristate
flabel metal2 s 439106 -960 439218 480 0 FreeSans 448 90 0 0 la_data_out[88]
port 385 nsew signal tristate
flabel metal2 s 442602 -960 442714 480 0 FreeSans 448 90 0 0 la_data_out[89]
port 386 nsew signal tristate
flabel metal2 s 155378 -960 155490 480 0 FreeSans 448 90 0 0 la_data_out[8]
port 387 nsew signal tristate
flabel metal2 s 446190 -960 446302 480 0 FreeSans 448 90 0 0 la_data_out[90]
port 388 nsew signal tristate
flabel metal2 s 449778 -960 449890 480 0 FreeSans 448 90 0 0 la_data_out[91]
port 389 nsew signal tristate
flabel metal2 s 453274 -960 453386 480 0 FreeSans 448 90 0 0 la_data_out[92]
port 390 nsew signal tristate
flabel metal2 s 456862 -960 456974 480 0 FreeSans 448 90 0 0 la_data_out[93]
port 391 nsew signal tristate
flabel metal2 s 460358 -960 460470 480 0 FreeSans 448 90 0 0 la_data_out[94]
port 392 nsew signal tristate
flabel metal2 s 463946 -960 464058 480 0 FreeSans 448 90 0 0 la_data_out[95]
port 393 nsew signal tristate
flabel metal2 s 467442 -960 467554 480 0 FreeSans 448 90 0 0 la_data_out[96]
port 394 nsew signal tristate
flabel metal2 s 471030 -960 471142 480 0 FreeSans 448 90 0 0 la_data_out[97]
port 395 nsew signal tristate
flabel metal2 s 474526 -960 474638 480 0 FreeSans 448 90 0 0 la_data_out[98]
port 396 nsew signal tristate
flabel metal2 s 478114 -960 478226 480 0 FreeSans 448 90 0 0 la_data_out[99]
port 397 nsew signal tristate
flabel metal2 s 158874 -960 158986 480 0 FreeSans 448 90 0 0 la_data_out[9]
port 398 nsew signal tristate
flabel metal2 s 128146 -960 128258 480 0 FreeSans 448 90 0 0 la_oenb[0]
port 399 nsew signal input
flabel metal2 s 482806 -960 482918 480 0 FreeSans 448 90 0 0 la_oenb[100]
port 400 nsew signal input
flabel metal2 s 486394 -960 486506 480 0 FreeSans 448 90 0 0 la_oenb[101]
port 401 nsew signal input
flabel metal2 s 489890 -960 490002 480 0 FreeSans 448 90 0 0 la_oenb[102]
port 402 nsew signal input
flabel metal2 s 493478 -960 493590 480 0 FreeSans 448 90 0 0 la_oenb[103]
port 403 nsew signal input
flabel metal2 s 497066 -960 497178 480 0 FreeSans 448 90 0 0 la_oenb[104]
port 404 nsew signal input
flabel metal2 s 500562 -960 500674 480 0 FreeSans 448 90 0 0 la_oenb[105]
port 405 nsew signal input
flabel metal2 s 504150 -960 504262 480 0 FreeSans 448 90 0 0 la_oenb[106]
port 406 nsew signal input
flabel metal2 s 507646 -960 507758 480 0 FreeSans 448 90 0 0 la_oenb[107]
port 407 nsew signal input
flabel metal2 s 511234 -960 511346 480 0 FreeSans 448 90 0 0 la_oenb[108]
port 408 nsew signal input
flabel metal2 s 514730 -960 514842 480 0 FreeSans 448 90 0 0 la_oenb[109]
port 409 nsew signal input
flabel metal2 s 163658 -960 163770 480 0 FreeSans 448 90 0 0 la_oenb[10]
port 410 nsew signal input
flabel metal2 s 518318 -960 518430 480 0 FreeSans 448 90 0 0 la_oenb[110]
port 411 nsew signal input
flabel metal2 s 521814 -960 521926 480 0 FreeSans 448 90 0 0 la_oenb[111]
port 412 nsew signal input
flabel metal2 s 525402 -960 525514 480 0 FreeSans 448 90 0 0 la_oenb[112]
port 413 nsew signal input
flabel metal2 s 528990 -960 529102 480 0 FreeSans 448 90 0 0 la_oenb[113]
port 414 nsew signal input
flabel metal2 s 532486 -960 532598 480 0 FreeSans 448 90 0 0 la_oenb[114]
port 415 nsew signal input
flabel metal2 s 536074 -960 536186 480 0 FreeSans 448 90 0 0 la_oenb[115]
port 416 nsew signal input
flabel metal2 s 539570 -960 539682 480 0 FreeSans 448 90 0 0 la_oenb[116]
port 417 nsew signal input
flabel metal2 s 543158 -960 543270 480 0 FreeSans 448 90 0 0 la_oenb[117]
port 418 nsew signal input
flabel metal2 s 546654 -960 546766 480 0 FreeSans 448 90 0 0 la_oenb[118]
port 419 nsew signal input
flabel metal2 s 550242 -960 550354 480 0 FreeSans 448 90 0 0 la_oenb[119]
port 420 nsew signal input
flabel metal2 s 167154 -960 167266 480 0 FreeSans 448 90 0 0 la_oenb[11]
port 421 nsew signal input
flabel metal2 s 553738 -960 553850 480 0 FreeSans 448 90 0 0 la_oenb[120]
port 422 nsew signal input
flabel metal2 s 557326 -960 557438 480 0 FreeSans 448 90 0 0 la_oenb[121]
port 423 nsew signal input
flabel metal2 s 560822 -960 560934 480 0 FreeSans 448 90 0 0 la_oenb[122]
port 424 nsew signal input
flabel metal2 s 564410 -960 564522 480 0 FreeSans 448 90 0 0 la_oenb[123]
port 425 nsew signal input
flabel metal2 s 567998 -960 568110 480 0 FreeSans 448 90 0 0 la_oenb[124]
port 426 nsew signal input
flabel metal2 s 571494 -960 571606 480 0 FreeSans 448 90 0 0 la_oenb[125]
port 427 nsew signal input
flabel metal2 s 575082 -960 575194 480 0 FreeSans 448 90 0 0 la_oenb[126]
port 428 nsew signal input
flabel metal2 s 578578 -960 578690 480 0 FreeSans 448 90 0 0 la_oenb[127]
port 429 nsew signal input
flabel metal2 s 170742 -960 170854 480 0 FreeSans 448 90 0 0 la_oenb[12]
port 430 nsew signal input
flabel metal2 s 174238 -960 174350 480 0 FreeSans 448 90 0 0 la_oenb[13]
port 431 nsew signal input
flabel metal2 s 177826 -960 177938 480 0 FreeSans 448 90 0 0 la_oenb[14]
port 432 nsew signal input
flabel metal2 s 181414 -960 181526 480 0 FreeSans 448 90 0 0 la_oenb[15]
port 433 nsew signal input
flabel metal2 s 184910 -960 185022 480 0 FreeSans 448 90 0 0 la_oenb[16]
port 434 nsew signal input
flabel metal2 s 188498 -960 188610 480 0 FreeSans 448 90 0 0 la_oenb[17]
port 435 nsew signal input
flabel metal2 s 191994 -960 192106 480 0 FreeSans 448 90 0 0 la_oenb[18]
port 436 nsew signal input
flabel metal2 s 195582 -960 195694 480 0 FreeSans 448 90 0 0 la_oenb[19]
port 437 nsew signal input
flabel metal2 s 131734 -960 131846 480 0 FreeSans 448 90 0 0 la_oenb[1]
port 438 nsew signal input
flabel metal2 s 199078 -960 199190 480 0 FreeSans 448 90 0 0 la_oenb[20]
port 439 nsew signal input
flabel metal2 s 202666 -960 202778 480 0 FreeSans 448 90 0 0 la_oenb[21]
port 440 nsew signal input
flabel metal2 s 206162 -960 206274 480 0 FreeSans 448 90 0 0 la_oenb[22]
port 441 nsew signal input
flabel metal2 s 209750 -960 209862 480 0 FreeSans 448 90 0 0 la_oenb[23]
port 442 nsew signal input
flabel metal2 s 213338 -960 213450 480 0 FreeSans 448 90 0 0 la_oenb[24]
port 443 nsew signal input
flabel metal2 s 216834 -960 216946 480 0 FreeSans 448 90 0 0 la_oenb[25]
port 444 nsew signal input
flabel metal2 s 220422 -960 220534 480 0 FreeSans 448 90 0 0 la_oenb[26]
port 445 nsew signal input
flabel metal2 s 223918 -960 224030 480 0 FreeSans 448 90 0 0 la_oenb[27]
port 446 nsew signal input
flabel metal2 s 227506 -960 227618 480 0 FreeSans 448 90 0 0 la_oenb[28]
port 447 nsew signal input
flabel metal2 s 231002 -960 231114 480 0 FreeSans 448 90 0 0 la_oenb[29]
port 448 nsew signal input
flabel metal2 s 135230 -960 135342 480 0 FreeSans 448 90 0 0 la_oenb[2]
port 449 nsew signal input
flabel metal2 s 234590 -960 234702 480 0 FreeSans 448 90 0 0 la_oenb[30]
port 450 nsew signal input
flabel metal2 s 238086 -960 238198 480 0 FreeSans 448 90 0 0 la_oenb[31]
port 451 nsew signal input
flabel metal2 s 241674 -960 241786 480 0 FreeSans 448 90 0 0 la_oenb[32]
port 452 nsew signal input
flabel metal2 s 245170 -960 245282 480 0 FreeSans 448 90 0 0 la_oenb[33]
port 453 nsew signal input
flabel metal2 s 248758 -960 248870 480 0 FreeSans 448 90 0 0 la_oenb[34]
port 454 nsew signal input
flabel metal2 s 252346 -960 252458 480 0 FreeSans 448 90 0 0 la_oenb[35]
port 455 nsew signal input
flabel metal2 s 255842 -960 255954 480 0 FreeSans 448 90 0 0 la_oenb[36]
port 456 nsew signal input
flabel metal2 s 259430 -960 259542 480 0 FreeSans 448 90 0 0 la_oenb[37]
port 457 nsew signal input
flabel metal2 s 262926 -960 263038 480 0 FreeSans 448 90 0 0 la_oenb[38]
port 458 nsew signal input
flabel metal2 s 266514 -960 266626 480 0 FreeSans 448 90 0 0 la_oenb[39]
port 459 nsew signal input
flabel metal2 s 138818 -960 138930 480 0 FreeSans 448 90 0 0 la_oenb[3]
port 460 nsew signal input
flabel metal2 s 270010 -960 270122 480 0 FreeSans 448 90 0 0 la_oenb[40]
port 461 nsew signal input
flabel metal2 s 273598 -960 273710 480 0 FreeSans 448 90 0 0 la_oenb[41]
port 462 nsew signal input
flabel metal2 s 277094 -960 277206 480 0 FreeSans 448 90 0 0 la_oenb[42]
port 463 nsew signal input
flabel metal2 s 280682 -960 280794 480 0 FreeSans 448 90 0 0 la_oenb[43]
port 464 nsew signal input
flabel metal2 s 284270 -960 284382 480 0 FreeSans 448 90 0 0 la_oenb[44]
port 465 nsew signal input
flabel metal2 s 287766 -960 287878 480 0 FreeSans 448 90 0 0 la_oenb[45]
port 466 nsew signal input
flabel metal2 s 291354 -960 291466 480 0 FreeSans 448 90 0 0 la_oenb[46]
port 467 nsew signal input
flabel metal2 s 294850 -960 294962 480 0 FreeSans 448 90 0 0 la_oenb[47]
port 468 nsew signal input
flabel metal2 s 298438 -960 298550 480 0 FreeSans 448 90 0 0 la_oenb[48]
port 469 nsew signal input
flabel metal2 s 301934 -960 302046 480 0 FreeSans 448 90 0 0 la_oenb[49]
port 470 nsew signal input
flabel metal2 s 142406 -960 142518 480 0 FreeSans 448 90 0 0 la_oenb[4]
port 471 nsew signal input
flabel metal2 s 305522 -960 305634 480 0 FreeSans 448 90 0 0 la_oenb[50]
port 472 nsew signal input
flabel metal2 s 309018 -960 309130 480 0 FreeSans 448 90 0 0 la_oenb[51]
port 473 nsew signal input
flabel metal2 s 312606 -960 312718 480 0 FreeSans 448 90 0 0 la_oenb[52]
port 474 nsew signal input
flabel metal2 s 316194 -960 316306 480 0 FreeSans 448 90 0 0 la_oenb[53]
port 475 nsew signal input
flabel metal2 s 319690 -960 319802 480 0 FreeSans 448 90 0 0 la_oenb[54]
port 476 nsew signal input
flabel metal2 s 323278 -960 323390 480 0 FreeSans 448 90 0 0 la_oenb[55]
port 477 nsew signal input
flabel metal2 s 326774 -960 326886 480 0 FreeSans 448 90 0 0 la_oenb[56]
port 478 nsew signal input
flabel metal2 s 330362 -960 330474 480 0 FreeSans 448 90 0 0 la_oenb[57]
port 479 nsew signal input
flabel metal2 s 333858 -960 333970 480 0 FreeSans 448 90 0 0 la_oenb[58]
port 480 nsew signal input
flabel metal2 s 337446 -960 337558 480 0 FreeSans 448 90 0 0 la_oenb[59]
port 481 nsew signal input
flabel metal2 s 145902 -960 146014 480 0 FreeSans 448 90 0 0 la_oenb[5]
port 482 nsew signal input
flabel metal2 s 340942 -960 341054 480 0 FreeSans 448 90 0 0 la_oenb[60]
port 483 nsew signal input
flabel metal2 s 344530 -960 344642 480 0 FreeSans 448 90 0 0 la_oenb[61]
port 484 nsew signal input
flabel metal2 s 348026 -960 348138 480 0 FreeSans 448 90 0 0 la_oenb[62]
port 485 nsew signal input
flabel metal2 s 351614 -960 351726 480 0 FreeSans 448 90 0 0 la_oenb[63]
port 486 nsew signal input
flabel metal2 s 355202 -960 355314 480 0 FreeSans 448 90 0 0 la_oenb[64]
port 487 nsew signal input
flabel metal2 s 358698 -960 358810 480 0 FreeSans 448 90 0 0 la_oenb[65]
port 488 nsew signal input
flabel metal2 s 362286 -960 362398 480 0 FreeSans 448 90 0 0 la_oenb[66]
port 489 nsew signal input
flabel metal2 s 365782 -960 365894 480 0 FreeSans 448 90 0 0 la_oenb[67]
port 490 nsew signal input
flabel metal2 s 369370 -960 369482 480 0 FreeSans 448 90 0 0 la_oenb[68]
port 491 nsew signal input
flabel metal2 s 372866 -960 372978 480 0 FreeSans 448 90 0 0 la_oenb[69]
port 492 nsew signal input
flabel metal2 s 149490 -960 149602 480 0 FreeSans 448 90 0 0 la_oenb[6]
port 493 nsew signal input
flabel metal2 s 376454 -960 376566 480 0 FreeSans 448 90 0 0 la_oenb[70]
port 494 nsew signal input
flabel metal2 s 379950 -960 380062 480 0 FreeSans 448 90 0 0 la_oenb[71]
port 495 nsew signal input
flabel metal2 s 383538 -960 383650 480 0 FreeSans 448 90 0 0 la_oenb[72]
port 496 nsew signal input
flabel metal2 s 387126 -960 387238 480 0 FreeSans 448 90 0 0 la_oenb[73]
port 497 nsew signal input
flabel metal2 s 390622 -960 390734 480 0 FreeSans 448 90 0 0 la_oenb[74]
port 498 nsew signal input
flabel metal2 s 394210 -960 394322 480 0 FreeSans 448 90 0 0 la_oenb[75]
port 499 nsew signal input
flabel metal2 s 397706 -960 397818 480 0 FreeSans 448 90 0 0 la_oenb[76]
port 500 nsew signal input
flabel metal2 s 401294 -960 401406 480 0 FreeSans 448 90 0 0 la_oenb[77]
port 501 nsew signal input
flabel metal2 s 404790 -960 404902 480 0 FreeSans 448 90 0 0 la_oenb[78]
port 502 nsew signal input
flabel metal2 s 408378 -960 408490 480 0 FreeSans 448 90 0 0 la_oenb[79]
port 503 nsew signal input
flabel metal2 s 152986 -960 153098 480 0 FreeSans 448 90 0 0 la_oenb[7]
port 504 nsew signal input
flabel metal2 s 411874 -960 411986 480 0 FreeSans 448 90 0 0 la_oenb[80]
port 505 nsew signal input
flabel metal2 s 415462 -960 415574 480 0 FreeSans 448 90 0 0 la_oenb[81]
port 506 nsew signal input
flabel metal2 s 418958 -960 419070 480 0 FreeSans 448 90 0 0 la_oenb[82]
port 507 nsew signal input
flabel metal2 s 422546 -960 422658 480 0 FreeSans 448 90 0 0 la_oenb[83]
port 508 nsew signal input
flabel metal2 s 426134 -960 426246 480 0 FreeSans 448 90 0 0 la_oenb[84]
port 509 nsew signal input
flabel metal2 s 429630 -960 429742 480 0 FreeSans 448 90 0 0 la_oenb[85]
port 510 nsew signal input
flabel metal2 s 433218 -960 433330 480 0 FreeSans 448 90 0 0 la_oenb[86]
port 511 nsew signal input
flabel metal2 s 436714 -960 436826 480 0 FreeSans 448 90 0 0 la_oenb[87]
port 512 nsew signal input
flabel metal2 s 440302 -960 440414 480 0 FreeSans 448 90 0 0 la_oenb[88]
port 513 nsew signal input
flabel metal2 s 443798 -960 443910 480 0 FreeSans 448 90 0 0 la_oenb[89]
port 514 nsew signal input
flabel metal2 s 156574 -960 156686 480 0 FreeSans 448 90 0 0 la_oenb[8]
port 515 nsew signal input
flabel metal2 s 447386 -960 447498 480 0 FreeSans 448 90 0 0 la_oenb[90]
port 516 nsew signal input
flabel metal2 s 450882 -960 450994 480 0 FreeSans 448 90 0 0 la_oenb[91]
port 517 nsew signal input
flabel metal2 s 454470 -960 454582 480 0 FreeSans 448 90 0 0 la_oenb[92]
port 518 nsew signal input
flabel metal2 s 458058 -960 458170 480 0 FreeSans 448 90 0 0 la_oenb[93]
port 519 nsew signal input
flabel metal2 s 461554 -960 461666 480 0 FreeSans 448 90 0 0 la_oenb[94]
port 520 nsew signal input
flabel metal2 s 465142 -960 465254 480 0 FreeSans 448 90 0 0 la_oenb[95]
port 521 nsew signal input
flabel metal2 s 468638 -960 468750 480 0 FreeSans 448 90 0 0 la_oenb[96]
port 522 nsew signal input
flabel metal2 s 472226 -960 472338 480 0 FreeSans 448 90 0 0 la_oenb[97]
port 523 nsew signal input
flabel metal2 s 475722 -960 475834 480 0 FreeSans 448 90 0 0 la_oenb[98]
port 524 nsew signal input
flabel metal2 s 479310 -960 479422 480 0 FreeSans 448 90 0 0 la_oenb[99]
port 525 nsew signal input
flabel metal2 s 160070 -960 160182 480 0 FreeSans 448 90 0 0 la_oenb[9]
port 526 nsew signal input
flabel metal2 s 579774 -960 579886 480 0 FreeSans 448 90 0 0 user_clock2
port 527 nsew signal input
flabel metal2 s 580970 -960 581082 480 0 FreeSans 448 90 0 0 user_irq[0]
port 528 nsew signal tristate
flabel metal2 s 582166 -960 582278 480 0 FreeSans 448 90 0 0 user_irq[1]
port 529 nsew signal tristate
flabel metal2 s 583362 -960 583474 480 0 FreeSans 448 90 0 0 user_irq[2]
port 530 nsew signal tristate
flabel metal4 s -2006 -934 -1386 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 -934 585930 -314 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 704250 585930 704870 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 585310 -934 585930 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 1794 -7654 2414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 37794 -7654 38414 12559 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 37794 677977 38414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 73794 -7654 74414 12559 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 73794 677977 74414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 109794 -7654 110414 12559 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 109794 677977 110414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 145794 -7654 146414 12559 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 145794 677977 146414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181794 -7654 182414 12559 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181794 677977 182414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 217794 -7654 218414 12559 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 217794 677977 218414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 253794 -7654 254414 12559 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 253794 677977 254414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 289794 -7654 290414 12559 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 289794 677977 290414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 325794 -7654 326414 12559 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 325794 677977 326414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 361794 -7654 362414 12559 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 361794 677977 362414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 397794 -7654 398414 12559 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 397794 677977 398414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 433794 -7654 434414 12559 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 433794 677977 434414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 469794 -7654 470414 12559 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 469794 677977 470414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 505794 -7654 506414 12559 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 505794 677977 506414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 541794 -7654 542414 12559 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 541794 677977 542414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 577794 -7654 578414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 2866 592650 3486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 38866 592650 39486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 74866 592650 75486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 110866 592650 111486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 146866 592650 147486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 182866 592650 183486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 218866 592650 219486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 254866 592650 255486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 290866 592650 291486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 326866 592650 327486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 362866 592650 363486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 398866 592650 399486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 434866 592650 435486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 470866 592650 471486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 506866 592650 507486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 542866 592650 543486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 578866 592650 579486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 614866 592650 615486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 650866 592650 651486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 686866 592650 687486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s -3926 -2854 -3306 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 -2854 587850 -2234 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 706170 587850 706790 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 587230 -2854 587850 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 9234 -7654 9854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 45234 -7654 45854 12559 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 45234 677977 45854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 81234 -7654 81854 12559 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 81234 677977 81854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 117234 -7654 117854 12559 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 117234 677977 117854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 153234 -7654 153854 12559 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 153234 677977 153854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 189234 -7654 189854 12559 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 189234 677977 189854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 225234 -7654 225854 12559 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 225234 677977 225854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 261234 -7654 261854 12559 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 261234 677977 261854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 297234 -7654 297854 12559 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 297234 677977 297854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 333234 -7654 333854 12559 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 333234 677977 333854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 369234 -7654 369854 12068 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 369234 678332 369854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 405234 -7654 405854 12559 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 405234 677977 405854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 441234 -7654 441854 12559 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 441234 677977 441854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 477234 -7654 477854 12068 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 477234 678332 477854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 513234 -7654 513854 12559 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 513234 677977 513854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 549234 -7654 549854 12559 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 549234 677977 549854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 10306 592650 10926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 46306 592650 46926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 82306 592650 82926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 118306 592650 118926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 154306 592650 154926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 190306 592650 190926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 226306 592650 226926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 262306 592650 262926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 298306 592650 298926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 334306 592650 334926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 370306 592650 370926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 406306 592650 406926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 442306 592650 442926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 478306 592650 478926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 514306 592650 514926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 550306 592650 550926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 586306 592650 586926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 622306 592650 622926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 658306 592650 658926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 694306 592650 694926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s -5846 -4774 -5226 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 -4774 589770 -4154 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 708090 589770 708710 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 589150 -4774 589770 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 17746 592650 18366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 53746 592650 54366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 89746 592650 90366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 125746 592650 126366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 161746 592650 162366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 197746 592650 198366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 233746 592650 234366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 269746 592650 270366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 305746 592650 306366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 341746 592650 342366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 377746 592650 378366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 413746 592650 414366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 449746 592650 450366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 485746 592650 486366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 521746 592650 522366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 557746 592650 558366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 593746 592650 594366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 629746 592650 630366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 665746 592650 666366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s -7766 -6694 -7146 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 -6694 591690 -6074 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 710010 591690 710630 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 591070 -6694 591690 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 25186 592650 25806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 61186 592650 61806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 97186 592650 97806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 133186 592650 133806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 169186 592650 169806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 205186 592650 205806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 241186 592650 241806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 277186 592650 277806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 313186 592650 313806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 349186 592650 349806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 385186 592650 385806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 421186 592650 421806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 457186 592650 457806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 493186 592650 493806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 529186 592650 529806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 565186 592650 565806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 601186 592650 601806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 637186 592650 637806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 673186 592650 673806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s -6806 -5734 -6186 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 -5734 590730 -5114 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 709050 590730 709670 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 590110 -5734 590730 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 21466 592650 22086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 57466 592650 58086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 93466 592650 94086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 129466 592650 130086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 165466 592650 166086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 201466 592650 202086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 237466 592650 238086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 273466 592650 274086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 309466 592650 310086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 345466 592650 346086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 381466 592650 382086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 417466 592650 418086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 453466 592650 454086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 489466 592650 490086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 525466 592650 526086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 561466 592650 562086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 597466 592650 598086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 633466 592650 634086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 669466 592650 670086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s -8726 -7654 -8106 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 -7654 592650 -7034 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 710970 592650 711590 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 592030 -7654 592650 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 567834 -7654 568454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 28906 592650 29526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 64906 592650 65526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 100906 592650 101526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 136906 592650 137526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 172906 592650 173526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 208906 592650 209526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 244906 592650 245526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 280906 592650 281526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 316906 592650 317526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 352906 592650 353526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 388906 592650 389526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 424906 592650 425526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 460906 592650 461526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 496906 592650 497526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 532906 592650 533526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 568906 592650 569526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 604906 592650 605526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 640906 592650 641526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 676906 592650 677526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s -2966 -1894 -2346 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 -1894 586890 -1274 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 705210 586890 705830 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 586270 -1894 586890 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 5514 -7654 6134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 41514 -7654 42134 12559 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 41514 677977 42134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 77514 -7654 78134 12068 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 77514 678332 78134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 113514 -7654 114134 12559 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 113514 677977 114134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 149514 -7654 150134 12559 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 149514 677977 150134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 185514 -7654 186134 12068 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 185514 678332 186134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 221514 -7654 222134 12559 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 221514 677977 222134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 257514 -7654 258134 12559 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 257514 677977 258134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 293514 -7654 294134 12559 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 293514 677977 294134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 329514 -7654 330134 12559 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 329514 677977 330134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 365514 -7654 366134 12559 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 365514 677977 366134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 401514 -7654 402134 12559 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 401514 677977 402134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 437514 -7654 438134 12559 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 437514 677977 438134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 473514 -7654 474134 12559 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 473514 677977 474134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 509514 -7654 510134 12559 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 509514 677977 510134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 545514 -7654 546134 12559 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 545514 677977 546134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 581514 -7654 582134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 6586 592650 7206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 42586 592650 43206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 78586 592650 79206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 114586 592650 115206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 150586 592650 151206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 186586 592650 187206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 222586 592650 223206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 258586 592650 259206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 294586 592650 295206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 330586 592650 331206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 366586 592650 367206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 402586 592650 403206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 438586 592650 439206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 474586 592650 475206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 510586 592650 511206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 546586 592650 547206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 582586 592650 583206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 618586 592650 619206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 654586 592650 655206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 690586 592650 691206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s -4886 -3814 -4266 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 -3814 588810 -3194 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 707130 588810 707750 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 588190 -3814 588810 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 12954 677977 13574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 48954 677977 49574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 84954 677977 85574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 120954 677977 121574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 156954 677977 157574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 192954 677977 193574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 228954 677977 229574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 264954 677977 265574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 300954 677977 301574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 336954 677977 337574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 372954 677977 373574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 408954 677977 409574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 444954 677977 445574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 480954 677977 481574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 516954 677977 517574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 552954 677977 553574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 14026 592650 14646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 50026 592650 50646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 86026 592650 86646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 122026 592650 122646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 158026 592650 158646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 194026 592650 194646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 230026 592650 230646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 266026 592650 266646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 302026 592650 302646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 338026 592650 338646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 374026 592650 374646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 410026 592650 410646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 446026 592650 446646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 482026 592650 482646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 518026 592650 518646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 554026 592650 554646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 590026 592650 590646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 626026 592650 626646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 662026 592650 662646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 698026 592650 698646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal2 s 542 -960 654 480 0 FreeSans 448 90 0 0 wb_clk_i
port 539 nsew signal input
flabel metal2 s 1646 -960 1758 480 0 FreeSans 448 90 0 0 wb_rst_i
port 540 nsew signal input
flabel metal2 s 2842 -960 2954 480 0 FreeSans 448 90 0 0 wbs_ack_o
port 541 nsew signal tristate
flabel metal2 s 7626 -960 7738 480 0 FreeSans 448 90 0 0 wbs_adr_i[0]
port 542 nsew signal input
flabel metal2 s 47830 -960 47942 480 0 FreeSans 448 90 0 0 wbs_adr_i[10]
port 543 nsew signal input
flabel metal2 s 51326 -960 51438 480 0 FreeSans 448 90 0 0 wbs_adr_i[11]
port 544 nsew signal input
flabel metal2 s 54914 -960 55026 480 0 FreeSans 448 90 0 0 wbs_adr_i[12]
port 545 nsew signal input
flabel metal2 s 58410 -960 58522 480 0 FreeSans 448 90 0 0 wbs_adr_i[13]
port 546 nsew signal input
flabel metal2 s 61998 -960 62110 480 0 FreeSans 448 90 0 0 wbs_adr_i[14]
port 547 nsew signal input
flabel metal2 s 65494 -960 65606 480 0 FreeSans 448 90 0 0 wbs_adr_i[15]
port 548 nsew signal input
flabel metal2 s 69082 -960 69194 480 0 FreeSans 448 90 0 0 wbs_adr_i[16]
port 549 nsew signal input
flabel metal2 s 72578 -960 72690 480 0 FreeSans 448 90 0 0 wbs_adr_i[17]
port 550 nsew signal input
flabel metal2 s 76166 -960 76278 480 0 FreeSans 448 90 0 0 wbs_adr_i[18]
port 551 nsew signal input
flabel metal2 s 79662 -960 79774 480 0 FreeSans 448 90 0 0 wbs_adr_i[19]
port 552 nsew signal input
flabel metal2 s 12318 -960 12430 480 0 FreeSans 448 90 0 0 wbs_adr_i[1]
port 553 nsew signal input
flabel metal2 s 83250 -960 83362 480 0 FreeSans 448 90 0 0 wbs_adr_i[20]
port 554 nsew signal input
flabel metal2 s 86838 -960 86950 480 0 FreeSans 448 90 0 0 wbs_adr_i[21]
port 555 nsew signal input
flabel metal2 s 90334 -960 90446 480 0 FreeSans 448 90 0 0 wbs_adr_i[22]
port 556 nsew signal input
flabel metal2 s 93922 -960 94034 480 0 FreeSans 448 90 0 0 wbs_adr_i[23]
port 557 nsew signal input
flabel metal2 s 97418 -960 97530 480 0 FreeSans 448 90 0 0 wbs_adr_i[24]
port 558 nsew signal input
flabel metal2 s 101006 -960 101118 480 0 FreeSans 448 90 0 0 wbs_adr_i[25]
port 559 nsew signal input
flabel metal2 s 104502 -960 104614 480 0 FreeSans 448 90 0 0 wbs_adr_i[26]
port 560 nsew signal input
flabel metal2 s 108090 -960 108202 480 0 FreeSans 448 90 0 0 wbs_adr_i[27]
port 561 nsew signal input
flabel metal2 s 111586 -960 111698 480 0 FreeSans 448 90 0 0 wbs_adr_i[28]
port 562 nsew signal input
flabel metal2 s 115174 -960 115286 480 0 FreeSans 448 90 0 0 wbs_adr_i[29]
port 563 nsew signal input
flabel metal2 s 17010 -960 17122 480 0 FreeSans 448 90 0 0 wbs_adr_i[2]
port 564 nsew signal input
flabel metal2 s 118762 -960 118874 480 0 FreeSans 448 90 0 0 wbs_adr_i[30]
port 565 nsew signal input
flabel metal2 s 122258 -960 122370 480 0 FreeSans 448 90 0 0 wbs_adr_i[31]
port 566 nsew signal input
flabel metal2 s 21794 -960 21906 480 0 FreeSans 448 90 0 0 wbs_adr_i[3]
port 567 nsew signal input
flabel metal2 s 26486 -960 26598 480 0 FreeSans 448 90 0 0 wbs_adr_i[4]
port 568 nsew signal input
flabel metal2 s 30074 -960 30186 480 0 FreeSans 448 90 0 0 wbs_adr_i[5]
port 569 nsew signal input
flabel metal2 s 33570 -960 33682 480 0 FreeSans 448 90 0 0 wbs_adr_i[6]
port 570 nsew signal input
flabel metal2 s 37158 -960 37270 480 0 FreeSans 448 90 0 0 wbs_adr_i[7]
port 571 nsew signal input
flabel metal2 s 40654 -960 40766 480 0 FreeSans 448 90 0 0 wbs_adr_i[8]
port 572 nsew signal input
flabel metal2 s 44242 -960 44354 480 0 FreeSans 448 90 0 0 wbs_adr_i[9]
port 573 nsew signal input
flabel metal2 s 4038 -960 4150 480 0 FreeSans 448 90 0 0 wbs_cyc_i
port 574 nsew signal input
flabel metal2 s 8730 -960 8842 480 0 FreeSans 448 90 0 0 wbs_dat_i[0]
port 575 nsew signal input
flabel metal2 s 48934 -960 49046 480 0 FreeSans 448 90 0 0 wbs_dat_i[10]
port 576 nsew signal input
flabel metal2 s 52522 -960 52634 480 0 FreeSans 448 90 0 0 wbs_dat_i[11]
port 577 nsew signal input
flabel metal2 s 56018 -960 56130 480 0 FreeSans 448 90 0 0 wbs_dat_i[12]
port 578 nsew signal input
flabel metal2 s 59606 -960 59718 480 0 FreeSans 448 90 0 0 wbs_dat_i[13]
port 579 nsew signal input
flabel metal2 s 63194 -960 63306 480 0 FreeSans 448 90 0 0 wbs_dat_i[14]
port 580 nsew signal input
flabel metal2 s 66690 -960 66802 480 0 FreeSans 448 90 0 0 wbs_dat_i[15]
port 581 nsew signal input
flabel metal2 s 70278 -960 70390 480 0 FreeSans 448 90 0 0 wbs_dat_i[16]
port 582 nsew signal input
flabel metal2 s 73774 -960 73886 480 0 FreeSans 448 90 0 0 wbs_dat_i[17]
port 583 nsew signal input
flabel metal2 s 77362 -960 77474 480 0 FreeSans 448 90 0 0 wbs_dat_i[18]
port 584 nsew signal input
flabel metal2 s 80858 -960 80970 480 0 FreeSans 448 90 0 0 wbs_dat_i[19]
port 585 nsew signal input
flabel metal2 s 13514 -960 13626 480 0 FreeSans 448 90 0 0 wbs_dat_i[1]
port 586 nsew signal input
flabel metal2 s 84446 -960 84558 480 0 FreeSans 448 90 0 0 wbs_dat_i[20]
port 587 nsew signal input
flabel metal2 s 87942 -960 88054 480 0 FreeSans 448 90 0 0 wbs_dat_i[21]
port 588 nsew signal input
flabel metal2 s 91530 -960 91642 480 0 FreeSans 448 90 0 0 wbs_dat_i[22]
port 589 nsew signal input
flabel metal2 s 95118 -960 95230 480 0 FreeSans 448 90 0 0 wbs_dat_i[23]
port 590 nsew signal input
flabel metal2 s 98614 -960 98726 480 0 FreeSans 448 90 0 0 wbs_dat_i[24]
port 591 nsew signal input
flabel metal2 s 102202 -960 102314 480 0 FreeSans 448 90 0 0 wbs_dat_i[25]
port 592 nsew signal input
flabel metal2 s 105698 -960 105810 480 0 FreeSans 448 90 0 0 wbs_dat_i[26]
port 593 nsew signal input
flabel metal2 s 109286 -960 109398 480 0 FreeSans 448 90 0 0 wbs_dat_i[27]
port 594 nsew signal input
flabel metal2 s 112782 -960 112894 480 0 FreeSans 448 90 0 0 wbs_dat_i[28]
port 595 nsew signal input
flabel metal2 s 116370 -960 116482 480 0 FreeSans 448 90 0 0 wbs_dat_i[29]
port 596 nsew signal input
flabel metal2 s 18206 -960 18318 480 0 FreeSans 448 90 0 0 wbs_dat_i[2]
port 597 nsew signal input
flabel metal2 s 119866 -960 119978 480 0 FreeSans 448 90 0 0 wbs_dat_i[30]
port 598 nsew signal input
flabel metal2 s 123454 -960 123566 480 0 FreeSans 448 90 0 0 wbs_dat_i[31]
port 599 nsew signal input
flabel metal2 s 22990 -960 23102 480 0 FreeSans 448 90 0 0 wbs_dat_i[3]
port 600 nsew signal input
flabel metal2 s 27682 -960 27794 480 0 FreeSans 448 90 0 0 wbs_dat_i[4]
port 601 nsew signal input
flabel metal2 s 31270 -960 31382 480 0 FreeSans 448 90 0 0 wbs_dat_i[5]
port 602 nsew signal input
flabel metal2 s 34766 -960 34878 480 0 FreeSans 448 90 0 0 wbs_dat_i[6]
port 603 nsew signal input
flabel metal2 s 38354 -960 38466 480 0 FreeSans 448 90 0 0 wbs_dat_i[7]
port 604 nsew signal input
flabel metal2 s 41850 -960 41962 480 0 FreeSans 448 90 0 0 wbs_dat_i[8]
port 605 nsew signal input
flabel metal2 s 45438 -960 45550 480 0 FreeSans 448 90 0 0 wbs_dat_i[9]
port 606 nsew signal input
flabel metal2 s 9926 -960 10038 480 0 FreeSans 448 90 0 0 wbs_dat_o[0]
port 607 nsew signal tristate
flabel metal2 s 50130 -960 50242 480 0 FreeSans 448 90 0 0 wbs_dat_o[10]
port 608 nsew signal tristate
flabel metal2 s 53718 -960 53830 480 0 FreeSans 448 90 0 0 wbs_dat_o[11]
port 609 nsew signal tristate
flabel metal2 s 57214 -960 57326 480 0 FreeSans 448 90 0 0 wbs_dat_o[12]
port 610 nsew signal tristate
flabel metal2 s 60802 -960 60914 480 0 FreeSans 448 90 0 0 wbs_dat_o[13]
port 611 nsew signal tristate
flabel metal2 s 64298 -960 64410 480 0 FreeSans 448 90 0 0 wbs_dat_o[14]
port 612 nsew signal tristate
flabel metal2 s 67886 -960 67998 480 0 FreeSans 448 90 0 0 wbs_dat_o[15]
port 613 nsew signal tristate
flabel metal2 s 71474 -960 71586 480 0 FreeSans 448 90 0 0 wbs_dat_o[16]
port 614 nsew signal tristate
flabel metal2 s 74970 -960 75082 480 0 FreeSans 448 90 0 0 wbs_dat_o[17]
port 615 nsew signal tristate
flabel metal2 s 78558 -960 78670 480 0 FreeSans 448 90 0 0 wbs_dat_o[18]
port 616 nsew signal tristate
flabel metal2 s 82054 -960 82166 480 0 FreeSans 448 90 0 0 wbs_dat_o[19]
port 617 nsew signal tristate
flabel metal2 s 14710 -960 14822 480 0 FreeSans 448 90 0 0 wbs_dat_o[1]
port 618 nsew signal tristate
flabel metal2 s 85642 -960 85754 480 0 FreeSans 448 90 0 0 wbs_dat_o[20]
port 619 nsew signal tristate
flabel metal2 s 89138 -960 89250 480 0 FreeSans 448 90 0 0 wbs_dat_o[21]
port 620 nsew signal tristate
flabel metal2 s 92726 -960 92838 480 0 FreeSans 448 90 0 0 wbs_dat_o[22]
port 621 nsew signal tristate
flabel metal2 s 96222 -960 96334 480 0 FreeSans 448 90 0 0 wbs_dat_o[23]
port 622 nsew signal tristate
flabel metal2 s 99810 -960 99922 480 0 FreeSans 448 90 0 0 wbs_dat_o[24]
port 623 nsew signal tristate
flabel metal2 s 103306 -960 103418 480 0 FreeSans 448 90 0 0 wbs_dat_o[25]
port 624 nsew signal tristate
flabel metal2 s 106894 -960 107006 480 0 FreeSans 448 90 0 0 wbs_dat_o[26]
port 625 nsew signal tristate
flabel metal2 s 110482 -960 110594 480 0 FreeSans 448 90 0 0 wbs_dat_o[27]
port 626 nsew signal tristate
flabel metal2 s 113978 -960 114090 480 0 FreeSans 448 90 0 0 wbs_dat_o[28]
port 627 nsew signal tristate
flabel metal2 s 117566 -960 117678 480 0 FreeSans 448 90 0 0 wbs_dat_o[29]
port 628 nsew signal tristate
flabel metal2 s 19402 -960 19514 480 0 FreeSans 448 90 0 0 wbs_dat_o[2]
port 629 nsew signal tristate
flabel metal2 s 121062 -960 121174 480 0 FreeSans 448 90 0 0 wbs_dat_o[30]
port 630 nsew signal tristate
flabel metal2 s 124650 -960 124762 480 0 FreeSans 448 90 0 0 wbs_dat_o[31]
port 631 nsew signal tristate
flabel metal2 s 24186 -960 24298 480 0 FreeSans 448 90 0 0 wbs_dat_o[3]
port 632 nsew signal tristate
flabel metal2 s 28878 -960 28990 480 0 FreeSans 448 90 0 0 wbs_dat_o[4]
port 633 nsew signal tristate
flabel metal2 s 32374 -960 32486 480 0 FreeSans 448 90 0 0 wbs_dat_o[5]
port 634 nsew signal tristate
flabel metal2 s 35962 -960 36074 480 0 FreeSans 448 90 0 0 wbs_dat_o[6]
port 635 nsew signal tristate
flabel metal2 s 39550 -960 39662 480 0 FreeSans 448 90 0 0 wbs_dat_o[7]
port 636 nsew signal tristate
flabel metal2 s 43046 -960 43158 480 0 FreeSans 448 90 0 0 wbs_dat_o[8]
port 637 nsew signal tristate
flabel metal2 s 46634 -960 46746 480 0 FreeSans 448 90 0 0 wbs_dat_o[9]
port 638 nsew signal tristate
flabel metal2 s 11122 -960 11234 480 0 FreeSans 448 90 0 0 wbs_sel_i[0]
port 639 nsew signal input
flabel metal2 s 15906 -960 16018 480 0 FreeSans 448 90 0 0 wbs_sel_i[1]
port 640 nsew signal input
flabel metal2 s 20598 -960 20710 480 0 FreeSans 448 90 0 0 wbs_sel_i[2]
port 641 nsew signal input
flabel metal2 s 25290 -960 25402 480 0 FreeSans 448 90 0 0 wbs_sel_i[3]
port 642 nsew signal input
flabel metal2 s 5234 -960 5346 480 0 FreeSans 448 90 0 0 wbs_stb_i
port 643 nsew signal input
flabel metal2 s 6430 -960 6542 480 0 FreeSans 448 90 0 0 wbs_we_i
port 644 nsew signal input
rlabel via4 538608 651336 538608 651336 0 vccd1
rlabel metal5 291962 694616 291962 694616 0 vccd2
rlabel metal5 291962 666056 291962 666056 0 vdda1
rlabel metal5 291962 673496 291962 673496 0 vdda2
rlabel metal5 291962 669776 291962 669776 0 vssa1
rlabel metal5 291962 677216 291962 677216 0 vssa2
rlabel via4 553968 655056 553968 655056 0 vssd1
rlabel metal5 291962 698336 291962 698336 0 vssd2
rlabel metal2 580198 284869 580198 284869 0 analog_io[0]
rlabel metal2 446154 701940 446154 701940 0 analog_io[10]
rlabel metal2 373398 678708 373398 678708 0 analog_io[11]
rlabel metal2 312034 678708 312034 678708 0 analog_io[12]
rlabel metal2 250486 678708 250486 678708 0 analog_io[13]
rlabel metal2 189168 678708 189168 678708 0 analog_io[14]
rlabel metal2 121670 701634 121670 701634 0 analog_io[15]
rlabel metal2 56626 682043 56626 682043 0 analog_io[16]
rlabel metal3 1878 697340 1878 697340 0 analog_io[17]
rlabel metal3 1924 645116 1924 645116 0 analog_io[18]
rlabel metal3 1556 593028 1556 593028 0 analog_io[19]
rlabel metal2 580198 338351 580198 338351 0 analog_io[1]
rlabel metal3 1878 540804 1878 540804 0 analog_io[20]
rlabel metal3 1878 488716 1878 488716 0 analog_io[21]
rlabel metal3 1648 436628 1648 436628 0 analog_io[22]
rlabel metal3 1878 384404 1878 384404 0 analog_io[23]
rlabel metal3 1694 332316 1694 332316 0 analog_io[24]
rlabel metal3 1878 280092 1878 280092 0 analog_io[25]
rlabel metal3 1878 228004 1878 228004 0 analog_io[26]
rlabel metal3 1878 175916 1878 175916 0 analog_io[27]
rlabel metal3 2200 123692 2200 123692 0 analog_io[28]
rlabel metal3 581218 391748 581218 391748 0 analog_io[2]
rlabel metal3 581954 444788 581954 444788 0 analog_io[3]
rlabel metal1 578726 496842 578726 496842 0 analog_io[4]
rlabel metal2 580198 550885 580198 550885 0 analog_io[5]
rlabel metal2 580198 603653 580198 603653 0 analog_io[6]
rlabel metal2 580198 657135 580198 657135 0 analog_io[7]
rlabel metal2 557766 678708 557766 678708 0 analog_io[8]
rlabel metal2 496310 678708 496310 678708 0 analog_io[9]
rlabel metal3 581218 6596 581218 6596 0 io_in[0]
rlabel metal3 581908 458116 581908 458116 0 io_in[10]
rlabel metal2 580198 510969 580198 510969 0 io_in[11]
rlabel metal2 579830 563703 579830 563703 0 io_in[12]
rlabel metal2 580198 617185 580198 617185 0 io_in[13]
rlabel via2 580198 670701 580198 670701 0 io_in[14]
rlabel metal2 542494 678708 542494 678708 0 io_in[15]
rlabel metal2 480946 678708 480946 678708 0 io_in[16]
rlabel metal2 429870 701940 429870 701940 0 io_in[17]
rlabel metal2 364366 691567 364366 691567 0 io_in[18]
rlabel metal2 296762 678708 296762 678708 0 io_in[19]
rlabel metal2 580198 46597 580198 46597 0 io_in[1]
rlabel metal2 235122 678708 235122 678708 0 io_in[20]
rlabel metal2 173666 678708 173666 678708 0 io_in[21]
rlabel metal2 112256 678708 112256 678708 0 io_in[22]
rlabel metal2 40204 703596 40204 703596 0 io_in[23]
rlabel metal3 1924 684284 1924 684284 0 io_in[24]
rlabel metal3 1970 632060 1970 632060 0 io_in[25]
rlabel metal3 1648 579972 1648 579972 0 io_in[26]
rlabel metal3 1878 527884 1878 527884 0 io_in[27]
rlabel metal3 1878 475660 1878 475660 0 io_in[28]
rlabel metal3 1878 423572 1878 423572 0 io_in[29]
rlabel metal2 580198 86547 580198 86547 0 io_in[2]
rlabel metal3 1878 371348 1878 371348 0 io_in[30]
rlabel metal3 1878 319260 1878 319260 0 io_in[31]
rlabel metal3 1694 267172 1694 267172 0 io_in[32]
rlabel metal3 1878 214948 1878 214948 0 io_in[33]
rlabel metal3 1924 162860 1924 162860 0 io_in[34]
rlabel metal3 1556 110636 1556 110636 0 io_in[35]
rlabel metal3 1878 71604 1878 71604 0 io_in[36]
rlabel metal3 1556 32436 1556 32436 0 io_in[37]
rlabel metal1 578956 126922 578956 126922 0 io_in[3]
rlabel metal2 577990 168368 577990 168368 0 io_in[4]
rlabel metal2 579554 206363 579554 206363 0 io_in[5]
rlabel metal2 580198 245225 580198 245225 0 io_in[6]
rlabel metal3 581954 298724 581954 298724 0 io_in[7]
rlabel metal2 579554 349129 579554 349129 0 io_in[8]
rlabel metal2 580198 404651 580198 404651 0 io_in[9]
rlabel metal3 581218 33116 581218 33116 0 io_oeb[0]
rlabel metal1 579140 484398 579140 484398 0 io_oeb[10]
rlabel metal2 580198 537319 580198 537319 0 io_oeb[11]
rlabel metal2 579830 590835 579830 590835 0 io_oeb[12]
rlabel metal2 580198 643569 580198 643569 0 io_oeb[13]
rlabel metal2 580198 697085 580198 697085 0 io_oeb[14]
rlabel metal2 527206 701940 527206 701940 0 io_oeb[15]
rlabel metal2 450218 678708 450218 678708 0 io_oeb[16]
rlabel metal2 388762 678708 388762 678708 0 io_oeb[17]
rlabel metal2 327306 678708 327306 678708 0 io_oeb[18]
rlabel metal2 265850 678708 265850 678708 0 io_oeb[19]
rlabel metal3 581218 72964 581218 72964 0 io_oeb[1]
rlabel metal2 204440 678708 204440 678708 0 io_oeb[20]
rlabel metal1 138966 699686 138966 699686 0 io_oeb[21]
rlabel metal2 81574 678708 81574 678708 0 io_oeb[22]
rlabel metal2 20072 678708 20072 678708 0 io_oeb[23]
rlabel metal3 1878 658172 1878 658172 0 io_oeb[24]
rlabel metal3 1924 606084 1924 606084 0 io_oeb[25]
rlabel metal3 1924 553860 1924 553860 0 io_oeb[26]
rlabel metal3 1694 501772 1694 501772 0 io_oeb[27]
rlabel metal3 1556 449548 1556 449548 0 io_oeb[28]
rlabel metal3 1878 397460 1878 397460 0 io_oeb[29]
rlabel metal3 581218 112812 581218 112812 0 io_oeb[2]
rlabel metal3 2200 345372 2200 345372 0 io_oeb[30]
rlabel metal3 1878 293148 1878 293148 0 io_oeb[31]
rlabel metal3 1878 241060 1878 241060 0 io_oeb[32]
rlabel metal3 1878 188836 1878 188836 0 io_oeb[33]
rlabel metal3 1786 136748 1786 136748 0 io_oeb[34]
rlabel metal3 1556 84660 1556 84660 0 io_oeb[35]
rlabel metal3 1556 45492 1556 45492 0 io_oeb[36]
rlabel metal3 1878 6460 1878 6460 0 io_oeb[37]
rlabel metal2 579554 155023 579554 155023 0 io_oeb[3]
rlabel metal2 579554 193545 579554 193545 0 io_oeb[4]
rlabel metal2 580198 232441 580198 232441 0 io_oeb[5]
rlabel metal2 579830 272051 579830 272051 0 io_oeb[6]
rlabel metal2 580198 323391 580198 323391 0 io_oeb[7]
rlabel metal3 581218 378420 581218 378420 0 io_oeb[8]
rlabel metal2 580198 431103 580198 431103 0 io_oeb[9]
rlabel metal3 581264 19788 581264 19788 0 io_out[0]
rlabel metal2 580014 471019 580014 471019 0 io_out[10]
rlabel via2 580198 524467 580198 524467 0 io_out[11]
rlabel metal2 580198 577269 580198 577269 0 io_out[12]
rlabel metal2 580198 630751 580198 630751 0 io_out[13]
rlabel metal2 580198 683519 580198 683519 0 io_out[14]
rlabel metal2 527252 678851 527252 678851 0 io_out[15]
rlabel metal2 465582 678708 465582 678708 0 io_out[16]
rlabel metal2 404126 678708 404126 678708 0 io_out[17]
rlabel metal2 348818 701940 348818 701940 0 io_out[18]
rlabel metal2 281214 678708 281214 678708 0 io_out[19]
rlabel metal3 581218 59636 581218 59636 0 io_out[1]
rlabel metal2 218454 703596 218454 703596 0 io_out[20]
rlabel metal2 158348 678708 158348 678708 0 io_out[21]
rlabel metal2 96892 678708 96892 678708 0 io_out[22]
rlabel metal2 23828 703596 23828 703596 0 io_out[23]
rlabel metal3 1970 671228 1970 671228 0 io_out[24]
rlabel metal3 1878 619140 1878 619140 0 io_out[25]
rlabel metal3 1878 566916 1878 566916 0 io_out[26]
rlabel metal3 1878 514828 1878 514828 0 io_out[27]
rlabel metal3 1878 462604 1878 462604 0 io_out[28]
rlabel metal3 1740 410516 1740 410516 0 io_out[29]
rlabel metal3 581218 99484 581218 99484 0 io_out[2]
rlabel metal3 1556 358428 1556 358428 0 io_out[30]
rlabel metal3 1878 306204 1878 306204 0 io_out[31]
rlabel metal3 1878 254116 1878 254116 0 io_out[32]
rlabel metal3 1832 201892 1832 201892 0 io_out[33]
rlabel metal3 1878 149804 1878 149804 0 io_out[34]
rlabel metal3 1556 97580 1556 97580 0 io_out[35]
rlabel metal3 1740 58548 1740 58548 0 io_out[36]
rlabel metal3 1556 19380 1556 19380 0 io_out[37]
rlabel metal3 581218 139332 581218 139332 0 io_out[3]
rlabel metal1 578588 179350 578588 179350 0 io_out[4]
rlabel metal1 580037 219402 580037 219402 0 io_out[5]
rlabel metal1 579669 258094 579669 258094 0 io_out[6]
rlabel metal2 580198 311967 580198 311967 0 io_out[7]
rlabel metal1 578956 364718 578956 364718 0 io_out[8]
rlabel metal2 580198 418217 580198 418217 0 io_out[9]
rlabel metal2 133860 9452 133860 9452 0 la_data_in[0]
rlabel metal2 480562 2183 480562 2183 0 la_data_in[100]
rlabel metal2 484058 1894 484058 1894 0 la_data_in[101]
rlabel metal2 487646 1690 487646 1690 0 la_data_in[102]
rlabel metal2 488566 6596 488566 6596 0 la_data_in[103]
rlabel metal2 494730 1962 494730 1962 0 la_data_in[104]
rlabel metal2 482034 10659 482034 10659 0 la_data_in[105]
rlabel metal2 501814 2166 501814 2166 0 la_data_in[106]
rlabel metal2 505402 1894 505402 1894 0 la_data_in[107]
rlabel metal2 508898 1928 508898 1928 0 la_data_in[108]
rlabel metal2 507886 6154 507886 6154 0 la_data_in[109]
rlabel metal2 161322 1894 161322 1894 0 la_data_in[10]
rlabel metal2 515982 1928 515982 1928 0 la_data_in[110]
rlabel metal2 519570 1962 519570 1962 0 la_data_in[111]
rlabel metal2 523066 1894 523066 1894 0 la_data_in[112]
rlabel metal2 526654 1758 526654 1758 0 la_data_in[113]
rlabel metal2 525734 6426 525734 6426 0 la_data_in[114]
rlabel metal2 533738 1928 533738 1928 0 la_data_in[115]
rlabel metal2 518466 10829 518466 10829 0 la_data_in[116]
rlabel metal2 521594 10455 521594 10455 0 la_data_in[117]
rlabel metal2 544410 1962 544410 1962 0 la_data_in[118]
rlabel metal2 528310 10761 528310 10761 0 la_data_in[119]
rlabel metal2 164910 1792 164910 1792 0 la_data_in[11]
rlabel metal2 545790 6256 545790 6256 0 la_data_in[120]
rlabel metal2 554990 1962 554990 1962 0 la_data_in[121]
rlabel metal2 558578 1996 558578 1996 0 la_data_in[122]
rlabel metal2 562074 1758 562074 1758 0 la_data_in[123]
rlabel metal2 565662 1860 565662 1860 0 la_data_in[124]
rlabel metal2 568921 340 568921 340 0 la_data_in[125]
rlabel metal1 551724 3774 551724 3774 0 la_data_in[126]
rlabel metal2 576334 2098 576334 2098 0 la_data_in[127]
rlabel metal1 172960 9486 172960 9486 0 la_data_in[12]
rlabel metal2 171994 2030 171994 2030 0 la_data_in[13]
rlabel metal2 175490 1894 175490 1894 0 la_data_in[14]
rlabel metal2 179078 1928 179078 1928 0 la_data_in[15]
rlabel metal2 182574 1758 182574 1758 0 la_data_in[16]
rlabel metal2 186162 1826 186162 1826 0 la_data_in[17]
rlabel metal2 193446 12036 193446 12036 0 la_data_in[18]
rlabel metal1 194902 9418 194902 9418 0 la_data_in[19]
rlabel metal2 136620 9452 136620 9452 0 la_data_in[1]
rlabel metal2 196834 2200 196834 2200 0 la_data_in[20]
rlabel metal1 201756 9486 201756 9486 0 la_data_in[21]
rlabel metal1 205206 9554 205206 9554 0 la_data_in[22]
rlabel metal2 209898 10251 209898 10251 0 la_data_in[23]
rlabel metal1 212060 9146 212060 9146 0 la_data_in[24]
rlabel metal1 215602 9486 215602 9486 0 la_data_in[25]
rlabel metal2 218086 4342 218086 4342 0 la_data_in[26]
rlabel metal1 222318 9418 222318 9418 0 la_data_in[27]
rlabel metal1 225814 9418 225814 9418 0 la_data_in[28]
rlabel via1 229126 9641 229126 9641 0 la_data_in[29]
rlabel metal2 132986 1656 132986 1656 0 la_data_in[2]
rlabel metal1 232760 8398 232760 8398 0 la_data_in[30]
rlabel metal1 236072 9486 236072 9486 0 la_data_in[31]
rlabel metal2 239630 12036 239630 12036 0 la_data_in[32]
rlabel metal2 243080 12036 243080 12036 0 la_data_in[33]
rlabel metal2 246185 340 246185 340 0 la_data_in[34]
rlabel metal2 249948 12036 249948 12036 0 la_data_in[35]
rlabel metal2 253352 12036 253352 12036 0 la_data_in[36]
rlabel metal1 256864 9486 256864 9486 0 la_data_in[37]
rlabel metal2 260682 1962 260682 1962 0 la_data_in[38]
rlabel metal1 263810 9146 263810 9146 0 la_data_in[39]
rlabel metal2 136482 2200 136482 2200 0 la_data_in[3]
rlabel metal2 267766 4342 267766 4342 0 la_data_in[40]
rlabel metal1 270664 9486 270664 9486 0 la_data_in[41]
rlabel metal2 274850 1843 274850 1843 0 la_data_in[42]
rlabel metal2 276690 10217 276690 10217 0 la_data_in[43]
rlabel metal2 281743 340 281743 340 0 la_data_in[44]
rlabel metal1 284372 9418 284372 9418 0 la_data_in[45]
rlabel metal2 289018 1656 289018 1656 0 la_data_in[46]
rlabel metal2 292606 1928 292606 1928 0 la_data_in[47]
rlabel metal2 296102 1690 296102 1690 0 la_data_in[48]
rlabel metal2 296562 10183 296562 10183 0 la_data_in[49]
rlabel metal2 140070 2030 140070 2030 0 la_data_in[4]
rlabel metal2 303186 1894 303186 1894 0 la_data_in[50]
rlabel metal2 306774 2030 306774 2030 0 la_data_in[51]
rlabel metal2 310270 1826 310270 1826 0 la_data_in[52]
rlabel metal2 313858 1894 313858 1894 0 la_data_in[53]
rlabel metal1 313858 8874 313858 8874 0 la_data_in[54]
rlabel metal2 320942 1826 320942 1826 0 la_data_in[55]
rlabel metal2 324438 1758 324438 1758 0 la_data_in[56]
rlabel metal2 328026 2166 328026 2166 0 la_data_in[57]
rlabel metal2 331614 1758 331614 1758 0 la_data_in[58]
rlabel metal2 335110 1826 335110 1826 0 la_data_in[59]
rlabel metal2 143566 1826 143566 1826 0 la_data_in[5]
rlabel metal2 335202 5337 335202 5337 0 la_data_in[60]
rlabel metal2 342194 1622 342194 1622 0 la_data_in[61]
rlabel metal2 345782 2200 345782 2200 0 la_data_in[62]
rlabel metal2 349278 1894 349278 1894 0 la_data_in[63]
rlabel metal2 352866 1962 352866 1962 0 la_data_in[64]
rlabel metal1 350704 9418 350704 9418 0 la_data_in[65]
rlabel metal1 353694 9418 353694 9418 0 la_data_in[66]
rlabel metal2 363538 1792 363538 1792 0 la_data_in[67]
rlabel metal2 367034 2200 367034 2200 0 la_data_in[68]
rlabel metal2 370622 1996 370622 1996 0 la_data_in[69]
rlabel metal2 153518 12036 153518 12036 0 la_data_in[6]
rlabel metal1 367264 9486 367264 9486 0 la_data_in[70]
rlabel metal1 370300 9418 370300 9418 0 la_data_in[71]
rlabel metal1 372968 9486 372968 9486 0 la_data_in[72]
rlabel metal2 384790 2166 384790 2166 0 la_data_in[73]
rlabel metal2 388286 1962 388286 1962 0 la_data_in[74]
rlabel metal2 391874 1656 391874 1656 0 la_data_in[75]
rlabel metal1 386860 9486 386860 9486 0 la_data_in[76]
rlabel metal1 389804 9486 389804 9486 0 la_data_in[77]
rlabel metal2 392610 10285 392610 10285 0 la_data_in[78]
rlabel metal2 406042 1928 406042 1928 0 la_data_in[79]
rlabel metal1 156400 9486 156400 9486 0 la_data_in[7]
rlabel metal2 409630 2166 409630 2166 0 la_data_in[80]
rlabel metal2 403466 6256 403466 6256 0 la_data_in[81]
rlabel metal1 406364 9418 406364 9418 0 la_data_in[82]
rlabel metal1 410182 9486 410182 9486 0 la_data_in[83]
rlabel metal2 423798 1928 423798 1928 0 la_data_in[84]
rlabel metal2 427294 1826 427294 1826 0 la_data_in[85]
rlabel metal2 430882 2064 430882 2064 0 la_data_in[86]
rlabel metal2 422326 6154 422326 6154 0 la_data_in[87]
rlabel metal1 426742 9146 426742 9146 0 la_data_in[88]
rlabel metal1 429364 9282 429364 9282 0 la_data_in[89]
rlabel metal2 154238 1826 154238 1826 0 la_data_in[8]
rlabel metal2 445050 1894 445050 1894 0 la_data_in[90]
rlabel metal2 435666 10523 435666 10523 0 la_data_in[91]
rlabel metal2 438794 10659 438794 10659 0 la_data_in[92]
rlabel metal2 442290 10625 442290 10625 0 la_data_in[93]
rlabel metal2 445602 10795 445602 10795 0 la_data_in[94]
rlabel metal2 462806 4988 462806 4988 0 la_data_in[95]
rlabel metal2 466302 4512 466302 4512 0 la_data_in[96]
rlabel metal2 469890 1928 469890 1928 0 la_data_in[97]
rlabel metal2 473478 1962 473478 1962 0 la_data_in[98]
rlabel metal2 462162 10523 462162 10523 0 la_data_in[99]
rlabel metal2 157826 2234 157826 2234 0 la_data_in[9]
rlabel metal2 133998 5031 133998 5031 0 la_data_out[0]
rlabel metal2 481758 2064 481758 2064 0 la_data_out[100]
rlabel metal2 485254 1928 485254 1928 0 la_data_out[101]
rlabel metal2 488842 1758 488842 1758 0 la_data_out[102]
rlabel metal2 492338 1928 492338 1928 0 la_data_out[103]
rlabel metal2 495926 1690 495926 1690 0 la_data_out[104]
rlabel metal2 482954 10795 482954 10795 0 la_data_out[105]
rlabel metal2 503010 1928 503010 1928 0 la_data_out[106]
rlabel metal2 506506 1792 506506 1792 0 la_data_out[107]
rlabel metal2 506506 6222 506506 6222 0 la_data_out[108]
rlabel metal2 513590 1826 513590 1826 0 la_data_out[109]
rlabel metal2 162518 1826 162518 1826 0 la_data_out[10]
rlabel metal2 517178 1860 517178 1860 0 la_data_out[110]
rlabel metal2 520766 2234 520766 2234 0 la_data_out[111]
rlabel metal2 524262 1792 524262 1792 0 la_data_out[112]
rlabel metal2 527850 1928 527850 1928 0 la_data_out[113]
rlabel metal2 526470 6120 526470 6120 0 la_data_out[114]
rlabel metal2 516074 10795 516074 10795 0 la_data_out[115]
rlabel metal2 519570 10659 519570 10659 0 la_data_out[116]
rlabel metal2 522882 10727 522882 10727 0 la_data_out[117]
rlabel metal2 545514 1656 545514 1656 0 la_data_out[118]
rlabel metal2 549102 2098 549102 2098 0 la_data_out[119]
rlabel metal2 171320 12036 171320 12036 0 la_data_out[11]
rlabel metal2 552690 1894 552690 1894 0 la_data_out[120]
rlabel metal2 556285 204 556285 204 0 la_data_out[121]
rlabel metal2 559774 2200 559774 2200 0 la_data_out[122]
rlabel metal2 563270 2234 563270 2234 0 la_data_out[123]
rlabel metal2 566858 1792 566858 1792 0 la_data_out[124]
rlabel metal2 570354 1843 570354 1843 0 la_data_out[125]
rlabel metal1 552644 3910 552644 3910 0 la_data_out[126]
rlabel metal2 577438 2064 577438 2064 0 la_data_out[127]
rlabel metal2 174356 12036 174356 12036 0 la_data_out[12]
rlabel metal2 173190 1758 173190 1758 0 la_data_out[13]
rlabel metal2 176686 1826 176686 1826 0 la_data_out[14]
rlabel metal2 180274 1962 180274 1962 0 la_data_out[15]
rlabel metal2 183770 1928 183770 1928 0 la_data_out[16]
rlabel metal2 190916 12036 190916 12036 0 la_data_out[17]
rlabel metal2 190854 1894 190854 1894 0 la_data_out[18]
rlabel metal2 194442 1826 194442 1826 0 la_data_out[19]
rlabel metal2 138000 8364 138000 8364 0 la_data_out[1]
rlabel metal2 197938 4342 197938 4342 0 la_data_out[20]
rlabel metal1 202906 9146 202906 9146 0 la_data_out[21]
rlabel metal1 206356 9418 206356 9418 0 la_data_out[22]
rlabel metal2 211186 10217 211186 10217 0 la_data_out[23]
rlabel metal1 213210 9010 213210 9010 0 la_data_out[24]
rlabel metal1 216614 9418 216614 9418 0 la_data_out[25]
rlabel metal2 219282 4376 219282 4376 0 la_data_out[26]
rlabel metal1 223468 9486 223468 9486 0 la_data_out[27]
rlabel metal1 227056 9486 227056 9486 0 la_data_out[28]
rlabel metal1 230322 8466 230322 8466 0 la_data_out[29]
rlabel metal2 134182 1690 134182 1690 0 la_data_out[2]
rlabel metal2 233926 12036 233926 12036 0 la_data_out[30]
rlabel metal2 237222 9452 237222 9452 0 la_data_out[31]
rlabel metal2 240343 340 240343 340 0 la_data_out[32]
rlabel metal2 244214 9452 244214 9452 0 la_data_out[33]
rlabel metal2 247634 12036 247634 12036 0 la_data_out[34]
rlabel metal2 251160 9452 251160 9452 0 la_data_out[35]
rlabel metal2 254465 340 254465 340 0 la_data_out[36]
rlabel metal2 257922 10217 257922 10217 0 la_data_out[37]
rlabel metal2 261356 12036 261356 12036 0 la_data_out[38]
rlabel metal1 264960 9486 264960 9486 0 la_data_out[39]
rlabel metal2 137678 2234 137678 2234 0 la_data_out[3]
rlabel metal2 268870 4444 268870 4444 0 la_data_out[40]
rlabel metal1 271814 9554 271814 9554 0 la_data_out[41]
rlabel metal2 276046 1707 276046 1707 0 la_data_out[42]
rlabel metal1 278668 9486 278668 9486 0 la_data_out[43]
rlabel metal2 283130 1911 283130 1911 0 la_data_out[44]
rlabel metal2 286626 1690 286626 1690 0 la_data_out[45]
rlabel metal2 290214 1690 290214 1690 0 la_data_out[46]
rlabel metal2 293710 1758 293710 1758 0 la_data_out[47]
rlabel metal1 294952 9418 294952 9418 0 la_data_out[48]
rlabel metal2 300794 1758 300794 1758 0 la_data_out[49]
rlabel metal2 141266 2098 141266 2098 0 la_data_out[4]
rlabel metal2 304382 1860 304382 1860 0 la_data_out[50]
rlabel metal2 307970 2098 307970 2098 0 la_data_out[51]
rlabel metal2 311466 1894 311466 1894 0 la_data_out[52]
rlabel metal2 315054 1758 315054 1758 0 la_data_out[53]
rlabel metal1 315054 9486 315054 9486 0 la_data_out[54]
rlabel metal2 322138 1894 322138 1894 0 la_data_out[55]
rlabel metal2 325634 1928 325634 1928 0 la_data_out[56]
rlabel metal2 329222 1894 329222 1894 0 la_data_out[57]
rlabel metal2 332718 1928 332718 1928 0 la_data_out[58]
rlabel metal1 331660 9486 331660 9486 0 la_data_out[59]
rlabel metal2 144762 1690 144762 1690 0 la_data_out[5]
rlabel metal2 334098 9452 334098 9452 0 la_data_out[60]
rlabel metal2 343390 1826 343390 1826 0 la_data_out[61]
rlabel metal2 346978 2234 346978 2234 0 la_data_out[62]
rlabel metal2 350474 1826 350474 1826 0 la_data_out[63]
rlabel metal2 354062 1622 354062 1622 0 la_data_out[64]
rlabel metal1 350796 9486 350796 9486 0 la_data_out[65]
rlabel metal2 353970 10489 353970 10489 0 la_data_out[66]
rlabel metal2 364642 2234 364642 2234 0 la_data_out[67]
rlabel metal2 368230 2098 368230 2098 0 la_data_out[68]
rlabel metal2 371726 1690 371726 1690 0 la_data_out[69]
rlabel metal2 154760 12036 154760 12036 0 la_data_out[6]
rlabel metal1 367678 9418 367678 9418 0 la_data_out[70]
rlabel metal1 371358 9486 371358 9486 0 la_data_out[71]
rlabel metal2 373750 10557 373750 10557 0 la_data_out[72]
rlabel metal2 385986 1826 385986 1826 0 la_data_out[73]
rlabel metal2 389482 1894 389482 1894 0 la_data_out[74]
rlabel metal2 393070 1690 393070 1690 0 la_data_out[75]
rlabel metal1 388102 9350 388102 9350 0 la_data_out[76]
rlabel metal1 391138 9418 391138 9418 0 la_data_out[77]
rlabel metal2 403650 2098 403650 2098 0 la_data_out[78]
rlabel metal2 407238 1894 407238 1894 0 la_data_out[79]
rlabel metal2 151846 1928 151846 1928 0 la_data_out[7]
rlabel metal2 410826 2132 410826 2132 0 la_data_out[80]
rlabel metal1 404018 9282 404018 9282 0 la_data_out[81]
rlabel metal1 407192 9486 407192 9486 0 la_data_out[82]
rlabel metal1 411332 9554 411332 9554 0 la_data_out[83]
rlabel metal2 424994 1860 424994 1860 0 la_data_out[84]
rlabel metal2 428490 2098 428490 2098 0 la_data_out[85]
rlabel metal2 432078 1962 432078 1962 0 la_data_out[86]
rlabel metal2 423706 9452 423706 9452 0 la_data_out[87]
rlabel metal1 427340 9486 427340 9486 0 la_data_out[88]
rlabel metal2 442658 2064 442658 2064 0 la_data_out[89]
rlabel metal2 155434 2200 155434 2200 0 la_data_out[8]
rlabel metal2 446246 4852 446246 4852 0 la_data_out[90]
rlabel metal1 437736 9282 437736 9282 0 la_data_out[91]
rlabel metal2 440082 10591 440082 10591 0 la_data_out[92]
rlabel metal2 443394 10727 443394 10727 0 la_data_out[93]
rlabel metal2 446706 10421 446706 10421 0 la_data_out[94]
rlabel metal2 464002 1928 464002 1928 0 la_data_out[95]
rlabel metal2 467498 4546 467498 4546 0 la_data_out[96]
rlabel metal2 470534 6069 470534 6069 0 la_data_out[97]
rlabel metal2 459954 10251 459954 10251 0 la_data_out[98]
rlabel metal2 463266 10829 463266 10829 0 la_data_out[99]
rlabel metal2 158930 1996 158930 1996 0 la_data_out[9]
rlabel metal1 134872 9350 134872 9350 0 la_oenb[0]
rlabel metal2 482862 1928 482862 1928 0 la_oenb[100]
rlabel metal2 486450 1656 486450 1656 0 la_oenb[101]
rlabel metal2 487186 6086 487186 6086 0 la_oenb[102]
rlabel metal2 493534 1758 493534 1758 0 la_oenb[103]
rlabel metal2 480930 10591 480930 10591 0 la_oenb[104]
rlabel metal2 500618 1690 500618 1690 0 la_oenb[105]
rlabel metal2 504206 1826 504206 1826 0 la_oenb[106]
rlabel metal2 507702 1758 507702 1758 0 la_oenb[107]
rlabel metal2 506782 6290 506782 6290 0 la_oenb[108]
rlabel metal2 514786 1894 514786 1894 0 la_oenb[109]
rlabel metal2 163714 2064 163714 2064 0 la_oenb[10]
rlabel metal2 500802 10557 500802 10557 0 la_oenb[110]
rlabel metal2 521870 1928 521870 1928 0 la_oenb[111]
rlabel metal2 525458 1860 525458 1860 0 la_oenb[112]
rlabel metal2 524262 6494 524262 6494 0 la_oenb[113]
rlabel metal2 527942 6528 527942 6528 0 la_oenb[114]
rlabel metal2 517362 10591 517362 10591 0 la_oenb[115]
rlabel metal2 520674 10523 520674 10523 0 la_oenb[116]
rlabel metal2 523986 10557 523986 10557 0 la_oenb[117]
rlabel metal2 546710 1843 546710 1843 0 la_oenb[118]
rlabel metal2 545054 6426 545054 6426 0 la_oenb[119]
rlabel metal2 172615 11764 172615 11764 0 la_oenb[11]
rlabel metal2 553794 2047 553794 2047 0 la_oenb[120]
rlabel metal2 557382 1928 557382 1928 0 la_oenb[121]
rlabel metal2 560878 2166 560878 2166 0 la_oenb[122]
rlabel metal2 564466 1979 564466 1979 0 la_oenb[123]
rlabel metal2 546680 12036 546680 12036 0 la_oenb[124]
rlabel metal2 571550 1911 571550 1911 0 la_oenb[125]
rlabel metal2 575138 2132 575138 2132 0 la_oenb[126]
rlabel metal2 578634 2030 578634 2030 0 la_oenb[127]
rlabel metal2 175598 12036 175598 12036 0 la_oenb[12]
rlabel metal2 174294 1928 174294 1928 0 la_oenb[13]
rlabel metal2 177882 2200 177882 2200 0 la_oenb[14]
rlabel metal2 181470 1894 181470 1894 0 la_oenb[15]
rlabel metal2 184966 1792 184966 1792 0 la_oenb[16]
rlabel metal2 192204 12036 192204 12036 0 la_oenb[17]
rlabel metal1 193752 9486 193752 9486 0 la_oenb[18]
rlabel metal2 195638 1792 195638 1792 0 la_oenb[19]
rlabel metal2 139380 9452 139380 9452 0 la_oenb[1]
rlabel metal2 199134 4784 199134 4784 0 la_oenb[20]
rlabel metal2 202722 1826 202722 1826 0 la_oenb[21]
rlabel metal1 207460 9486 207460 9486 0 la_oenb[22]
rlabel metal1 210910 9486 210910 9486 0 la_oenb[23]
rlabel metal1 214360 9418 214360 9418 0 la_oenb[24]
rlabel metal1 217764 9486 217764 9486 0 la_oenb[25]
rlabel metal1 221352 9486 221352 9486 0 la_oenb[26]
rlabel metal1 224618 8738 224618 8738 0 la_oenb[27]
rlabel metal1 228068 9418 228068 9418 0 la_oenb[28]
rlabel metal1 231472 8738 231472 8738 0 la_oenb[29]
rlabel metal2 135286 1792 135286 1792 0 la_oenb[2]
rlabel metal2 235076 12036 235076 12036 0 la_oenb[30]
rlabel metal2 238142 4342 238142 4342 0 la_oenb[31]
rlabel metal2 241930 12036 241930 12036 0 la_oenb[32]
rlabel metal2 245334 12036 245334 12036 0 la_oenb[33]
rlabel metal2 248623 340 248623 340 0 la_oenb[34]
rlabel metal2 252248 12036 252248 12036 0 la_oenb[35]
rlabel metal2 255652 12036 255652 12036 0 la_oenb[36]
rlabel metal2 259486 1911 259486 1911 0 la_oenb[37]
rlabel metal1 262568 9486 262568 9486 0 la_oenb[38]
rlabel metal1 266110 8874 266110 8874 0 la_oenb[39]
rlabel metal2 138874 1996 138874 1996 0 la_oenb[3]
rlabel metal1 269514 9146 269514 9146 0 la_oenb[40]
rlabel metal1 272964 9418 272964 9418 0 la_oenb[41]
rlabel metal1 276368 9214 276368 9214 0 la_oenb[42]
rlabel metal2 280738 1690 280738 1690 0 la_oenb[43]
rlabel metal2 284326 1911 284326 1911 0 la_oenb[44]
rlabel metal2 287822 2098 287822 2098 0 la_oenb[45]
rlabel metal2 291410 1843 291410 1843 0 la_oenb[46]
rlabel metal2 294906 1928 294906 1928 0 la_oenb[47]
rlabel metal1 295780 9486 295780 9486 0 la_oenb[48]
rlabel metal2 301990 1928 301990 1928 0 la_oenb[49]
rlabel metal2 142462 1894 142462 1894 0 la_oenb[4]
rlabel metal2 305578 1962 305578 1962 0 la_oenb[50]
rlabel metal2 309074 1928 309074 1928 0 la_oenb[51]
rlabel metal2 312662 1928 312662 1928 0 la_oenb[52]
rlabel metal1 312524 9486 312524 9486 0 la_oenb[53]
rlabel metal2 315330 10285 315330 10285 0 la_oenb[54]
rlabel metal2 323334 1792 323334 1792 0 la_oenb[55]
rlabel metal2 326830 2234 326830 2234 0 la_oenb[56]
rlabel metal2 330418 1826 330418 1826 0 la_oenb[57]
rlabel metal2 333914 1894 333914 1894 0 la_oenb[58]
rlabel metal1 332902 9350 332902 9350 0 la_oenb[59]
rlabel metal2 152276 12036 152276 12036 0 la_oenb[5]
rlabel metal2 335202 10183 335202 10183 0 la_oenb[60]
rlabel metal2 344586 1792 344586 1792 0 la_oenb[61]
rlabel metal2 348082 1928 348082 1928 0 la_oenb[62]
rlabel metal2 351670 1860 351670 1860 0 la_oenb[63]
rlabel metal1 349462 8602 349462 8602 0 la_oenb[64]
rlabel metal1 352498 9486 352498 9486 0 la_oenb[65]
rlabel metal2 362342 1690 362342 1690 0 la_oenb[66]
rlabel metal2 365838 2166 365838 2166 0 la_oenb[67]
rlabel metal2 369426 2064 369426 2064 0 la_oenb[68]
rlabel metal2 372922 1894 372922 1894 0 la_oenb[69]
rlabel metal2 156055 11764 156055 11764 0 la_oenb[6]
rlabel metal1 369012 8602 369012 8602 0 la_oenb[70]
rlabel metal1 372140 9010 372140 9010 0 la_oenb[71]
rlabel metal2 383594 1656 383594 1656 0 la_oenb[72]
rlabel metal2 387182 2064 387182 2064 0 la_oenb[73]
rlabel metal2 390678 2030 390678 2030 0 la_oenb[74]
rlabel metal1 386768 3638 386768 3638 0 la_oenb[75]
rlabel metal1 389206 8874 389206 8874 0 la_oenb[76]
rlabel metal1 392012 9486 392012 9486 0 la_oenb[77]
rlabel metal2 404846 2030 404846 2030 0 la_oenb[78]
rlabel metal2 408434 2064 408434 2064 0 la_oenb[79]
rlabel metal2 153042 1622 153042 1622 0 la_oenb[7]
rlabel metal2 411930 1996 411930 1996 0 la_oenb[80]
rlabel metal1 405444 8738 405444 8738 0 la_oenb[81]
rlabel metal1 408296 9486 408296 9486 0 la_oenb[82]
rlabel metal2 422602 1996 422602 1996 0 la_oenb[83]
rlabel metal2 426190 2234 426190 2234 0 la_oenb[84]
rlabel metal2 429686 1894 429686 1894 0 la_oenb[85]
rlabel metal2 423062 6290 423062 6290 0 la_oenb[86]
rlabel metal1 425362 8602 425362 8602 0 la_oenb[87]
rlabel metal2 427570 10557 427570 10557 0 la_oenb[88]
rlabel metal2 443854 1962 443854 1962 0 la_oenb[89]
rlabel metal2 156630 1656 156630 1656 0 la_oenb[8]
rlabel metal2 434562 10489 434562 10489 0 la_oenb[90]
rlabel metal1 438380 9418 438380 9418 0 la_oenb[91]
rlabel metal2 441186 10319 441186 10319 0 la_oenb[92]
rlabel metal2 444314 10761 444314 10761 0 la_oenb[93]
rlabel metal2 461610 4682 461610 4682 0 la_oenb[94]
rlabel metal2 465198 1911 465198 1911 0 la_oenb[95]
rlabel metal2 468694 4444 468694 4444 0 la_oenb[96]
rlabel metal2 472282 1911 472282 1911 0 la_oenb[97]
rlabel metal2 475778 1928 475778 1928 0 la_oenb[98]
rlabel metal2 464370 10557 464370 10557 0 la_oenb[99]
rlabel metal2 160126 2030 160126 2030 0 la_oenb[9]
rlabel metal2 579830 1894 579830 1894 0 user_clock2
rlabel metal2 581026 1962 581026 1962 0 user_irq[0]
rlabel metal2 582222 2047 582222 2047 0 user_irq[1]
rlabel metal2 583418 1996 583418 1996 0 user_irq[2]
rlabel metal2 598 2064 598 2064 0 wb_clk_i
rlabel metal2 1702 1894 1702 1894 0 wb_rst_i
rlabel metal2 2898 2098 2898 2098 0 wbs_ack_o
rlabel metal2 18078 3706 18078 3706 0 wbs_adr_i[0]
rlabel metal2 60766 10625 60766 10625 0 wbs_adr_i[10]
rlabel metal1 61686 9418 61686 9418 0 wbs_adr_i[11]
rlabel metal2 60950 6460 60950 6460 0 wbs_adr_i[12]
rlabel metal2 58466 2234 58466 2234 0 wbs_adr_i[13]
rlabel metal2 62054 2200 62054 2200 0 wbs_adr_i[14]
rlabel metal2 77326 10625 77326 10625 0 wbs_adr_i[15]
rlabel metal1 78384 9486 78384 9486 0 wbs_adr_i[16]
rlabel metal2 79994 6460 79994 6460 0 wbs_adr_i[17]
rlabel metal2 76222 1690 76222 1690 0 wbs_adr_i[18]
rlabel metal2 79718 2234 79718 2234 0 wbs_adr_i[19]
rlabel metal2 12374 1962 12374 1962 0 wbs_adr_i[1]
rlabel metal2 83306 1928 83306 1928 0 wbs_adr_i[20]
rlabel metal2 97198 10591 97198 10591 0 wbs_adr_i[21]
rlabel metal1 98992 9010 98992 9010 0 wbs_adr_i[22]
rlabel metal2 93978 1622 93978 1622 0 wbs_adr_i[23]
rlabel metal2 97474 2234 97474 2234 0 wbs_adr_i[24]
rlabel metal2 101062 2132 101062 2132 0 wbs_adr_i[25]
rlabel metal2 113758 10183 113758 10183 0 wbs_adr_i[26]
rlabel metal1 115966 9486 115966 9486 0 wbs_adr_i[27]
rlabel metal1 119232 9010 119232 9010 0 wbs_adr_i[28]
rlabel metal2 115230 1860 115230 1860 0 wbs_adr_i[29]
rlabel metal2 17066 1758 17066 1758 0 wbs_adr_i[2]
rlabel metal2 118818 2166 118818 2166 0 wbs_adr_i[30]
rlabel metal2 122314 2098 122314 2098 0 wbs_adr_i[31]
rlabel metal2 21850 2098 21850 2098 0 wbs_adr_i[3]
rlabel metal2 40894 10727 40894 10727 0 wbs_adr_i[4]
rlabel metal1 40112 9554 40112 9554 0 wbs_adr_i[5]
rlabel metal2 41354 6494 41354 6494 0 wbs_adr_i[6]
rlabel metal2 37214 1928 37214 1928 0 wbs_adr_i[7]
rlabel metal2 40710 1826 40710 1826 0 wbs_adr_i[8]
rlabel metal2 44298 2132 44298 2132 0 wbs_adr_i[9]
rlabel metal2 4094 2132 4094 2132 0 wbs_cyc_i
rlabel metal1 21160 9486 21160 9486 0 wbs_dat_i[0]
rlabel metal1 58696 8874 58696 8874 0 wbs_dat_i[10]
rlabel metal2 60582 5916 60582 5916 0 wbs_dat_i[11]
rlabel metal2 56074 1656 56074 1656 0 wbs_dat_i[12]
rlabel metal2 59662 1962 59662 1962 0 wbs_dat_i[13]
rlabel metal2 63250 1996 63250 1996 0 wbs_dat_i[14]
rlabel metal2 78706 10523 78706 10523 0 wbs_dat_i[15]
rlabel metal1 78844 9622 78844 9622 0 wbs_dat_i[16]
rlabel metal2 80546 6018 80546 6018 0 wbs_dat_i[17]
rlabel metal2 77418 2200 77418 2200 0 wbs_dat_i[18]
rlabel metal2 80914 2098 80914 2098 0 wbs_dat_i[19]
rlabel metal2 23322 6324 23322 6324 0 wbs_dat_i[1]
rlabel metal2 95266 10183 95266 10183 0 wbs_dat_i[20]
rlabel metal1 96094 9486 96094 9486 0 wbs_dat_i[21]
rlabel metal1 100050 9486 100050 9486 0 wbs_dat_i[22]
rlabel metal2 95174 1894 95174 1894 0 wbs_dat_i[23]
rlabel metal2 98670 1758 98670 1758 0 wbs_dat_i[24]
rlabel metal2 102258 1894 102258 1894 0 wbs_dat_i[25]
rlabel metal2 114862 10591 114862 10591 0 wbs_dat_i[26]
rlabel metal1 117714 9418 117714 9418 0 wbs_dat_i[27]
rlabel metal1 120106 9418 120106 9418 0 wbs_dat_i[28]
rlabel metal2 116426 2234 116426 2234 0 wbs_dat_i[29]
rlabel metal2 18262 1928 18262 1928 0 wbs_dat_i[2]
rlabel metal2 119922 1894 119922 1894 0 wbs_dat_i[30]
rlabel metal2 123510 1690 123510 1690 0 wbs_dat_i[31]
rlabel metal2 23046 1996 23046 1996 0 wbs_dat_i[3]
rlabel metal2 41998 10761 41998 10761 0 wbs_dat_i[4]
rlabel metal2 37306 6426 37306 6426 0 wbs_dat_i[5]
rlabel metal2 41538 6460 41538 6460 0 wbs_dat_i[6]
rlabel metal2 38410 1690 38410 1690 0 wbs_dat_i[7]
rlabel metal2 41906 2030 41906 2030 0 wbs_dat_i[8]
rlabel metal2 45494 1894 45494 1894 0 wbs_dat_i[9]
rlabel metal1 23782 8874 23782 8874 0 wbs_dat_o[0]
rlabel metal1 59846 9282 59846 9282 0 wbs_dat_o[10]
rlabel metal2 60030 6188 60030 6188 0 wbs_dat_o[11]
rlabel metal2 57270 1928 57270 1928 0 wbs_dat_o[12]
rlabel metal2 60858 1894 60858 1894 0 wbs_dat_o[13]
rlabel metal2 64354 2064 64354 2064 0 wbs_dat_o[14]
rlabel metal1 77096 9418 77096 9418 0 wbs_dat_o[15]
rlabel metal1 80730 9554 80730 9554 0 wbs_dat_o[16]
rlabel metal2 75026 1928 75026 1928 0 wbs_dat_o[17]
rlabel metal2 78614 1826 78614 1826 0 wbs_dat_o[18]
rlabel metal2 82110 1962 82110 1962 0 wbs_dat_o[19]
rlabel metal2 24978 6732 24978 6732 0 wbs_dat_o[1]
rlabel metal2 96094 10625 96094 10625 0 wbs_dat_o[20]
rlabel metal2 95266 5507 95266 5507 0 wbs_dat_o[21]
rlabel metal1 101108 9418 101108 9418 0 wbs_dat_o[22]
rlabel metal2 96278 1860 96278 1860 0 wbs_dat_o[23]
rlabel metal2 99866 2064 99866 2064 0 wbs_dat_o[24]
rlabel metal2 103362 1928 103362 1928 0 wbs_dat_o[25]
rlabel metal1 114632 9418 114632 9418 0 wbs_dat_o[26]
rlabel metal1 118956 9486 118956 9486 0 wbs_dat_o[27]
rlabel metal2 114034 1690 114034 1690 0 wbs_dat_o[28]
rlabel metal2 117622 1826 117622 1826 0 wbs_dat_o[29]
rlabel metal2 19458 1894 19458 1894 0 wbs_dat_o[2]
rlabel metal2 121118 2030 121118 2030 0 wbs_dat_o[30]
rlabel metal2 132526 10848 132526 10848 0 wbs_dat_o[31]
rlabel metal2 24242 2166 24242 2166 0 wbs_dat_o[3]
rlabel metal2 43102 10693 43102 10693 0 wbs_dat_o[4]
rlabel metal2 39330 6018 39330 6018 0 wbs_dat_o[5]
rlabel metal2 36018 1656 36018 1656 0 wbs_dat_o[6]
rlabel metal2 39606 2234 39606 2234 0 wbs_dat_o[7]
rlabel metal2 43102 2064 43102 2064 0 wbs_dat_o[8]
rlabel metal2 59662 10489 59662 10489 0 wbs_dat_o[9]
rlabel metal2 11178 2030 11178 2030 0 wbs_sel_i[0]
rlabel metal2 23414 6426 23414 6426 0 wbs_sel_i[1]
rlabel metal2 20654 1826 20654 1826 0 wbs_sel_i[2]
rlabel metal2 25346 2064 25346 2064 0 wbs_sel_i[3]
rlabel metal2 5290 2234 5290 2234 0 wbs_stb_i
rlabel metal2 6486 1996 6486 1996 0 wbs_we_i
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
