magic
tech sky130A
magscale 1 2
timestamp 1669232171
<< obsli1 >>
rect 1104 2159 553012 664241
<< obsm1 >>
rect 382 2128 553012 664420
<< metal2 >>
rect 8206 665948 8262 666748
rect 23570 665948 23626 666748
rect 38934 665948 38990 666748
rect 54298 665948 54354 666748
rect 69662 665948 69718 666748
rect 85026 665948 85082 666748
rect 100390 665948 100446 666748
rect 115754 665948 115810 666748
rect 131118 665948 131174 666748
rect 146482 665948 146538 666748
rect 161846 665948 161902 666748
rect 177210 665948 177266 666748
rect 192574 665948 192630 666748
rect 207938 665948 207994 666748
rect 223302 665948 223358 666748
rect 238666 665948 238722 666748
rect 254030 665948 254086 666748
rect 269394 665948 269450 666748
rect 284758 665948 284814 666748
rect 300122 665948 300178 666748
rect 315486 665948 315542 666748
rect 330850 665948 330906 666748
rect 346214 665948 346270 666748
rect 361578 665948 361634 666748
rect 376942 665948 376998 666748
rect 392306 665948 392362 666748
rect 407670 665948 407726 666748
rect 423034 665948 423090 666748
rect 438398 665948 438454 666748
rect 453762 665948 453818 666748
rect 469126 665948 469182 666748
rect 484490 665948 484546 666748
rect 499854 665948 499910 666748
rect 515218 665948 515274 666748
rect 530582 665948 530638 666748
rect 545946 665948 546002 666748
rect 4894 0 4950 800
rect 5998 0 6054 800
rect 7102 0 7158 800
rect 8206 0 8262 800
rect 9310 0 9366 800
rect 10414 0 10470 800
rect 11518 0 11574 800
rect 12622 0 12678 800
rect 13726 0 13782 800
rect 14830 0 14886 800
rect 15934 0 15990 800
rect 17038 0 17094 800
rect 18142 0 18198 800
rect 19246 0 19302 800
rect 20350 0 20406 800
rect 21454 0 21510 800
rect 22558 0 22614 800
rect 23662 0 23718 800
rect 24766 0 24822 800
rect 25870 0 25926 800
rect 26974 0 27030 800
rect 28078 0 28134 800
rect 29182 0 29238 800
rect 30286 0 30342 800
rect 31390 0 31446 800
rect 32494 0 32550 800
rect 33598 0 33654 800
rect 34702 0 34758 800
rect 35806 0 35862 800
rect 36910 0 36966 800
rect 38014 0 38070 800
rect 39118 0 39174 800
rect 40222 0 40278 800
rect 41326 0 41382 800
rect 42430 0 42486 800
rect 43534 0 43590 800
rect 44638 0 44694 800
rect 45742 0 45798 800
rect 46846 0 46902 800
rect 47950 0 48006 800
rect 49054 0 49110 800
rect 50158 0 50214 800
rect 51262 0 51318 800
rect 52366 0 52422 800
rect 53470 0 53526 800
rect 54574 0 54630 800
rect 55678 0 55734 800
rect 56782 0 56838 800
rect 57886 0 57942 800
rect 58990 0 59046 800
rect 60094 0 60150 800
rect 61198 0 61254 800
rect 62302 0 62358 800
rect 63406 0 63462 800
rect 64510 0 64566 800
rect 65614 0 65670 800
rect 66718 0 66774 800
rect 67822 0 67878 800
rect 68926 0 68982 800
rect 70030 0 70086 800
rect 71134 0 71190 800
rect 72238 0 72294 800
rect 73342 0 73398 800
rect 74446 0 74502 800
rect 75550 0 75606 800
rect 76654 0 76710 800
rect 77758 0 77814 800
rect 78862 0 78918 800
rect 79966 0 80022 800
rect 81070 0 81126 800
rect 82174 0 82230 800
rect 83278 0 83334 800
rect 84382 0 84438 800
rect 85486 0 85542 800
rect 86590 0 86646 800
rect 87694 0 87750 800
rect 88798 0 88854 800
rect 89902 0 89958 800
rect 91006 0 91062 800
rect 92110 0 92166 800
rect 93214 0 93270 800
rect 94318 0 94374 800
rect 95422 0 95478 800
rect 96526 0 96582 800
rect 97630 0 97686 800
rect 98734 0 98790 800
rect 99838 0 99894 800
rect 100942 0 100998 800
rect 102046 0 102102 800
rect 103150 0 103206 800
rect 104254 0 104310 800
rect 105358 0 105414 800
rect 106462 0 106518 800
rect 107566 0 107622 800
rect 108670 0 108726 800
rect 109774 0 109830 800
rect 110878 0 110934 800
rect 111982 0 112038 800
rect 113086 0 113142 800
rect 114190 0 114246 800
rect 115294 0 115350 800
rect 116398 0 116454 800
rect 117502 0 117558 800
rect 118606 0 118662 800
rect 119710 0 119766 800
rect 120814 0 120870 800
rect 121918 0 121974 800
rect 123022 0 123078 800
rect 124126 0 124182 800
rect 125230 0 125286 800
rect 126334 0 126390 800
rect 127438 0 127494 800
rect 128542 0 128598 800
rect 129646 0 129702 800
rect 130750 0 130806 800
rect 131854 0 131910 800
rect 132958 0 133014 800
rect 134062 0 134118 800
rect 135166 0 135222 800
rect 136270 0 136326 800
rect 137374 0 137430 800
rect 138478 0 138534 800
rect 139582 0 139638 800
rect 140686 0 140742 800
rect 141790 0 141846 800
rect 142894 0 142950 800
rect 143998 0 144054 800
rect 145102 0 145158 800
rect 146206 0 146262 800
rect 147310 0 147366 800
rect 148414 0 148470 800
rect 149518 0 149574 800
rect 150622 0 150678 800
rect 151726 0 151782 800
rect 152830 0 152886 800
rect 153934 0 153990 800
rect 155038 0 155094 800
rect 156142 0 156198 800
rect 157246 0 157302 800
rect 158350 0 158406 800
rect 159454 0 159510 800
rect 160558 0 160614 800
rect 161662 0 161718 800
rect 162766 0 162822 800
rect 163870 0 163926 800
rect 164974 0 165030 800
rect 166078 0 166134 800
rect 167182 0 167238 800
rect 168286 0 168342 800
rect 169390 0 169446 800
rect 170494 0 170550 800
rect 171598 0 171654 800
rect 172702 0 172758 800
rect 173806 0 173862 800
rect 174910 0 174966 800
rect 176014 0 176070 800
rect 177118 0 177174 800
rect 178222 0 178278 800
rect 179326 0 179382 800
rect 180430 0 180486 800
rect 181534 0 181590 800
rect 182638 0 182694 800
rect 183742 0 183798 800
rect 184846 0 184902 800
rect 185950 0 186006 800
rect 187054 0 187110 800
rect 188158 0 188214 800
rect 189262 0 189318 800
rect 190366 0 190422 800
rect 191470 0 191526 800
rect 192574 0 192630 800
rect 193678 0 193734 800
rect 194782 0 194838 800
rect 195886 0 195942 800
rect 196990 0 197046 800
rect 198094 0 198150 800
rect 199198 0 199254 800
rect 200302 0 200358 800
rect 201406 0 201462 800
rect 202510 0 202566 800
rect 203614 0 203670 800
rect 204718 0 204774 800
rect 205822 0 205878 800
rect 206926 0 206982 800
rect 208030 0 208086 800
rect 209134 0 209190 800
rect 210238 0 210294 800
rect 211342 0 211398 800
rect 212446 0 212502 800
rect 213550 0 213606 800
rect 214654 0 214710 800
rect 215758 0 215814 800
rect 216862 0 216918 800
rect 217966 0 218022 800
rect 219070 0 219126 800
rect 220174 0 220230 800
rect 221278 0 221334 800
rect 222382 0 222438 800
rect 223486 0 223542 800
rect 224590 0 224646 800
rect 225694 0 225750 800
rect 226798 0 226854 800
rect 227902 0 227958 800
rect 229006 0 229062 800
rect 230110 0 230166 800
rect 231214 0 231270 800
rect 232318 0 232374 800
rect 233422 0 233478 800
rect 234526 0 234582 800
rect 235630 0 235686 800
rect 236734 0 236790 800
rect 237838 0 237894 800
rect 238942 0 238998 800
rect 240046 0 240102 800
rect 241150 0 241206 800
rect 242254 0 242310 800
rect 243358 0 243414 800
rect 244462 0 244518 800
rect 245566 0 245622 800
rect 246670 0 246726 800
rect 247774 0 247830 800
rect 248878 0 248934 800
rect 249982 0 250038 800
rect 251086 0 251142 800
rect 252190 0 252246 800
rect 253294 0 253350 800
rect 254398 0 254454 800
rect 255502 0 255558 800
rect 256606 0 256662 800
rect 257710 0 257766 800
rect 258814 0 258870 800
rect 259918 0 259974 800
rect 261022 0 261078 800
rect 262126 0 262182 800
rect 263230 0 263286 800
rect 264334 0 264390 800
rect 265438 0 265494 800
rect 266542 0 266598 800
rect 267646 0 267702 800
rect 268750 0 268806 800
rect 269854 0 269910 800
rect 270958 0 271014 800
rect 272062 0 272118 800
rect 273166 0 273222 800
rect 274270 0 274326 800
rect 275374 0 275430 800
rect 276478 0 276534 800
rect 277582 0 277638 800
rect 278686 0 278742 800
rect 279790 0 279846 800
rect 280894 0 280950 800
rect 281998 0 282054 800
rect 283102 0 283158 800
rect 284206 0 284262 800
rect 285310 0 285366 800
rect 286414 0 286470 800
rect 287518 0 287574 800
rect 288622 0 288678 800
rect 289726 0 289782 800
rect 290830 0 290886 800
rect 291934 0 291990 800
rect 293038 0 293094 800
rect 294142 0 294198 800
rect 295246 0 295302 800
rect 296350 0 296406 800
rect 297454 0 297510 800
rect 298558 0 298614 800
rect 299662 0 299718 800
rect 300766 0 300822 800
rect 301870 0 301926 800
rect 302974 0 303030 800
rect 304078 0 304134 800
rect 305182 0 305238 800
rect 306286 0 306342 800
rect 307390 0 307446 800
rect 308494 0 308550 800
rect 309598 0 309654 800
rect 310702 0 310758 800
rect 311806 0 311862 800
rect 312910 0 312966 800
rect 314014 0 314070 800
rect 315118 0 315174 800
rect 316222 0 316278 800
rect 317326 0 317382 800
rect 318430 0 318486 800
rect 319534 0 319590 800
rect 320638 0 320694 800
rect 321742 0 321798 800
rect 322846 0 322902 800
rect 323950 0 324006 800
rect 325054 0 325110 800
rect 326158 0 326214 800
rect 327262 0 327318 800
rect 328366 0 328422 800
rect 329470 0 329526 800
rect 330574 0 330630 800
rect 331678 0 331734 800
rect 332782 0 332838 800
rect 333886 0 333942 800
rect 334990 0 335046 800
rect 336094 0 336150 800
rect 337198 0 337254 800
rect 338302 0 338358 800
rect 339406 0 339462 800
rect 340510 0 340566 800
rect 341614 0 341670 800
rect 342718 0 342774 800
rect 343822 0 343878 800
rect 344926 0 344982 800
rect 346030 0 346086 800
rect 347134 0 347190 800
rect 348238 0 348294 800
rect 349342 0 349398 800
rect 350446 0 350502 800
rect 351550 0 351606 800
rect 352654 0 352710 800
rect 353758 0 353814 800
rect 354862 0 354918 800
rect 355966 0 356022 800
rect 357070 0 357126 800
rect 358174 0 358230 800
rect 359278 0 359334 800
rect 360382 0 360438 800
rect 361486 0 361542 800
rect 362590 0 362646 800
rect 363694 0 363750 800
rect 364798 0 364854 800
rect 365902 0 365958 800
rect 367006 0 367062 800
rect 368110 0 368166 800
rect 369214 0 369270 800
rect 370318 0 370374 800
rect 371422 0 371478 800
rect 372526 0 372582 800
rect 373630 0 373686 800
rect 374734 0 374790 800
rect 375838 0 375894 800
rect 376942 0 376998 800
rect 378046 0 378102 800
rect 379150 0 379206 800
rect 380254 0 380310 800
rect 381358 0 381414 800
rect 382462 0 382518 800
rect 383566 0 383622 800
rect 384670 0 384726 800
rect 385774 0 385830 800
rect 386878 0 386934 800
rect 387982 0 388038 800
rect 389086 0 389142 800
rect 390190 0 390246 800
rect 391294 0 391350 800
rect 392398 0 392454 800
rect 393502 0 393558 800
rect 394606 0 394662 800
rect 395710 0 395766 800
rect 396814 0 396870 800
rect 397918 0 397974 800
rect 399022 0 399078 800
rect 400126 0 400182 800
rect 401230 0 401286 800
rect 402334 0 402390 800
rect 403438 0 403494 800
rect 404542 0 404598 800
rect 405646 0 405702 800
rect 406750 0 406806 800
rect 407854 0 407910 800
rect 408958 0 409014 800
rect 410062 0 410118 800
rect 411166 0 411222 800
rect 412270 0 412326 800
rect 413374 0 413430 800
rect 414478 0 414534 800
rect 415582 0 415638 800
rect 416686 0 416742 800
rect 417790 0 417846 800
rect 418894 0 418950 800
rect 419998 0 420054 800
rect 421102 0 421158 800
rect 422206 0 422262 800
rect 423310 0 423366 800
rect 424414 0 424470 800
rect 425518 0 425574 800
rect 426622 0 426678 800
rect 427726 0 427782 800
rect 428830 0 428886 800
rect 429934 0 429990 800
rect 431038 0 431094 800
rect 432142 0 432198 800
rect 433246 0 433302 800
rect 434350 0 434406 800
rect 435454 0 435510 800
rect 436558 0 436614 800
rect 437662 0 437718 800
rect 438766 0 438822 800
rect 439870 0 439926 800
rect 440974 0 441030 800
rect 442078 0 442134 800
rect 443182 0 443238 800
rect 444286 0 444342 800
rect 445390 0 445446 800
rect 446494 0 446550 800
rect 447598 0 447654 800
rect 448702 0 448758 800
rect 449806 0 449862 800
rect 450910 0 450966 800
rect 452014 0 452070 800
rect 453118 0 453174 800
rect 454222 0 454278 800
rect 455326 0 455382 800
rect 456430 0 456486 800
rect 457534 0 457590 800
rect 458638 0 458694 800
rect 459742 0 459798 800
rect 460846 0 460902 800
rect 461950 0 462006 800
rect 463054 0 463110 800
rect 464158 0 464214 800
rect 465262 0 465318 800
rect 466366 0 466422 800
rect 467470 0 467526 800
rect 468574 0 468630 800
rect 469678 0 469734 800
rect 470782 0 470838 800
rect 471886 0 471942 800
rect 472990 0 473046 800
rect 474094 0 474150 800
rect 475198 0 475254 800
rect 476302 0 476358 800
rect 477406 0 477462 800
rect 478510 0 478566 800
rect 479614 0 479670 800
rect 480718 0 480774 800
rect 481822 0 481878 800
rect 482926 0 482982 800
rect 484030 0 484086 800
rect 485134 0 485190 800
rect 486238 0 486294 800
rect 487342 0 487398 800
rect 488446 0 488502 800
rect 489550 0 489606 800
rect 490654 0 490710 800
rect 491758 0 491814 800
rect 492862 0 492918 800
rect 493966 0 494022 800
rect 495070 0 495126 800
rect 496174 0 496230 800
rect 497278 0 497334 800
rect 498382 0 498438 800
rect 499486 0 499542 800
rect 500590 0 500646 800
rect 501694 0 501750 800
rect 502798 0 502854 800
rect 503902 0 503958 800
rect 505006 0 505062 800
rect 506110 0 506166 800
rect 507214 0 507270 800
rect 508318 0 508374 800
rect 509422 0 509478 800
rect 510526 0 510582 800
rect 511630 0 511686 800
rect 512734 0 512790 800
rect 513838 0 513894 800
rect 514942 0 514998 800
rect 516046 0 516102 800
rect 517150 0 517206 800
rect 518254 0 518310 800
rect 519358 0 519414 800
rect 520462 0 520518 800
rect 521566 0 521622 800
rect 522670 0 522726 800
rect 523774 0 523830 800
rect 524878 0 524934 800
rect 525982 0 526038 800
rect 527086 0 527142 800
rect 528190 0 528246 800
rect 529294 0 529350 800
rect 530398 0 530454 800
rect 531502 0 531558 800
rect 532606 0 532662 800
rect 533710 0 533766 800
rect 534814 0 534870 800
rect 535918 0 535974 800
rect 537022 0 537078 800
rect 538126 0 538182 800
rect 539230 0 539286 800
rect 540334 0 540390 800
rect 541438 0 541494 800
rect 542542 0 542598 800
rect 543646 0 543702 800
rect 544750 0 544806 800
rect 545854 0 545910 800
rect 546958 0 547014 800
rect 548062 0 548118 800
rect 549166 0 549222 800
<< obsm2 >>
rect 388 665892 8150 666074
rect 8318 665892 23514 666074
rect 23682 665892 38878 666074
rect 39046 665892 54242 666074
rect 54410 665892 69606 666074
rect 69774 665892 84970 666074
rect 85138 665892 100334 666074
rect 100502 665892 115698 666074
rect 115866 665892 131062 666074
rect 131230 665892 146426 666074
rect 146594 665892 161790 666074
rect 161958 665892 177154 666074
rect 177322 665892 192518 666074
rect 192686 665892 207882 666074
rect 208050 665892 223246 666074
rect 223414 665892 238610 666074
rect 238778 665892 253974 666074
rect 254142 665892 269338 666074
rect 269506 665892 284702 666074
rect 284870 665892 300066 666074
rect 300234 665892 315430 666074
rect 315598 665892 330794 666074
rect 330962 665892 346158 666074
rect 346326 665892 361522 666074
rect 361690 665892 376886 666074
rect 377054 665892 392250 666074
rect 392418 665892 407614 666074
rect 407782 665892 422978 666074
rect 423146 665892 438342 666074
rect 438510 665892 453706 666074
rect 453874 665892 469070 666074
rect 469238 665892 484434 666074
rect 484602 665892 499798 666074
rect 499966 665892 515162 666074
rect 515330 665892 530526 666074
rect 530694 665892 545890 666074
rect 546058 665892 552624 666074
rect 388 856 552624 665892
rect 388 734 4838 856
rect 5006 734 5942 856
rect 6110 734 7046 856
rect 7214 734 8150 856
rect 8318 734 9254 856
rect 9422 734 10358 856
rect 10526 734 11462 856
rect 11630 734 12566 856
rect 12734 734 13670 856
rect 13838 734 14774 856
rect 14942 734 15878 856
rect 16046 734 16982 856
rect 17150 734 18086 856
rect 18254 734 19190 856
rect 19358 734 20294 856
rect 20462 734 21398 856
rect 21566 734 22502 856
rect 22670 734 23606 856
rect 23774 734 24710 856
rect 24878 734 25814 856
rect 25982 734 26918 856
rect 27086 734 28022 856
rect 28190 734 29126 856
rect 29294 734 30230 856
rect 30398 734 31334 856
rect 31502 734 32438 856
rect 32606 734 33542 856
rect 33710 734 34646 856
rect 34814 734 35750 856
rect 35918 734 36854 856
rect 37022 734 37958 856
rect 38126 734 39062 856
rect 39230 734 40166 856
rect 40334 734 41270 856
rect 41438 734 42374 856
rect 42542 734 43478 856
rect 43646 734 44582 856
rect 44750 734 45686 856
rect 45854 734 46790 856
rect 46958 734 47894 856
rect 48062 734 48998 856
rect 49166 734 50102 856
rect 50270 734 51206 856
rect 51374 734 52310 856
rect 52478 734 53414 856
rect 53582 734 54518 856
rect 54686 734 55622 856
rect 55790 734 56726 856
rect 56894 734 57830 856
rect 57998 734 58934 856
rect 59102 734 60038 856
rect 60206 734 61142 856
rect 61310 734 62246 856
rect 62414 734 63350 856
rect 63518 734 64454 856
rect 64622 734 65558 856
rect 65726 734 66662 856
rect 66830 734 67766 856
rect 67934 734 68870 856
rect 69038 734 69974 856
rect 70142 734 71078 856
rect 71246 734 72182 856
rect 72350 734 73286 856
rect 73454 734 74390 856
rect 74558 734 75494 856
rect 75662 734 76598 856
rect 76766 734 77702 856
rect 77870 734 78806 856
rect 78974 734 79910 856
rect 80078 734 81014 856
rect 81182 734 82118 856
rect 82286 734 83222 856
rect 83390 734 84326 856
rect 84494 734 85430 856
rect 85598 734 86534 856
rect 86702 734 87638 856
rect 87806 734 88742 856
rect 88910 734 89846 856
rect 90014 734 90950 856
rect 91118 734 92054 856
rect 92222 734 93158 856
rect 93326 734 94262 856
rect 94430 734 95366 856
rect 95534 734 96470 856
rect 96638 734 97574 856
rect 97742 734 98678 856
rect 98846 734 99782 856
rect 99950 734 100886 856
rect 101054 734 101990 856
rect 102158 734 103094 856
rect 103262 734 104198 856
rect 104366 734 105302 856
rect 105470 734 106406 856
rect 106574 734 107510 856
rect 107678 734 108614 856
rect 108782 734 109718 856
rect 109886 734 110822 856
rect 110990 734 111926 856
rect 112094 734 113030 856
rect 113198 734 114134 856
rect 114302 734 115238 856
rect 115406 734 116342 856
rect 116510 734 117446 856
rect 117614 734 118550 856
rect 118718 734 119654 856
rect 119822 734 120758 856
rect 120926 734 121862 856
rect 122030 734 122966 856
rect 123134 734 124070 856
rect 124238 734 125174 856
rect 125342 734 126278 856
rect 126446 734 127382 856
rect 127550 734 128486 856
rect 128654 734 129590 856
rect 129758 734 130694 856
rect 130862 734 131798 856
rect 131966 734 132902 856
rect 133070 734 134006 856
rect 134174 734 135110 856
rect 135278 734 136214 856
rect 136382 734 137318 856
rect 137486 734 138422 856
rect 138590 734 139526 856
rect 139694 734 140630 856
rect 140798 734 141734 856
rect 141902 734 142838 856
rect 143006 734 143942 856
rect 144110 734 145046 856
rect 145214 734 146150 856
rect 146318 734 147254 856
rect 147422 734 148358 856
rect 148526 734 149462 856
rect 149630 734 150566 856
rect 150734 734 151670 856
rect 151838 734 152774 856
rect 152942 734 153878 856
rect 154046 734 154982 856
rect 155150 734 156086 856
rect 156254 734 157190 856
rect 157358 734 158294 856
rect 158462 734 159398 856
rect 159566 734 160502 856
rect 160670 734 161606 856
rect 161774 734 162710 856
rect 162878 734 163814 856
rect 163982 734 164918 856
rect 165086 734 166022 856
rect 166190 734 167126 856
rect 167294 734 168230 856
rect 168398 734 169334 856
rect 169502 734 170438 856
rect 170606 734 171542 856
rect 171710 734 172646 856
rect 172814 734 173750 856
rect 173918 734 174854 856
rect 175022 734 175958 856
rect 176126 734 177062 856
rect 177230 734 178166 856
rect 178334 734 179270 856
rect 179438 734 180374 856
rect 180542 734 181478 856
rect 181646 734 182582 856
rect 182750 734 183686 856
rect 183854 734 184790 856
rect 184958 734 185894 856
rect 186062 734 186998 856
rect 187166 734 188102 856
rect 188270 734 189206 856
rect 189374 734 190310 856
rect 190478 734 191414 856
rect 191582 734 192518 856
rect 192686 734 193622 856
rect 193790 734 194726 856
rect 194894 734 195830 856
rect 195998 734 196934 856
rect 197102 734 198038 856
rect 198206 734 199142 856
rect 199310 734 200246 856
rect 200414 734 201350 856
rect 201518 734 202454 856
rect 202622 734 203558 856
rect 203726 734 204662 856
rect 204830 734 205766 856
rect 205934 734 206870 856
rect 207038 734 207974 856
rect 208142 734 209078 856
rect 209246 734 210182 856
rect 210350 734 211286 856
rect 211454 734 212390 856
rect 212558 734 213494 856
rect 213662 734 214598 856
rect 214766 734 215702 856
rect 215870 734 216806 856
rect 216974 734 217910 856
rect 218078 734 219014 856
rect 219182 734 220118 856
rect 220286 734 221222 856
rect 221390 734 222326 856
rect 222494 734 223430 856
rect 223598 734 224534 856
rect 224702 734 225638 856
rect 225806 734 226742 856
rect 226910 734 227846 856
rect 228014 734 228950 856
rect 229118 734 230054 856
rect 230222 734 231158 856
rect 231326 734 232262 856
rect 232430 734 233366 856
rect 233534 734 234470 856
rect 234638 734 235574 856
rect 235742 734 236678 856
rect 236846 734 237782 856
rect 237950 734 238886 856
rect 239054 734 239990 856
rect 240158 734 241094 856
rect 241262 734 242198 856
rect 242366 734 243302 856
rect 243470 734 244406 856
rect 244574 734 245510 856
rect 245678 734 246614 856
rect 246782 734 247718 856
rect 247886 734 248822 856
rect 248990 734 249926 856
rect 250094 734 251030 856
rect 251198 734 252134 856
rect 252302 734 253238 856
rect 253406 734 254342 856
rect 254510 734 255446 856
rect 255614 734 256550 856
rect 256718 734 257654 856
rect 257822 734 258758 856
rect 258926 734 259862 856
rect 260030 734 260966 856
rect 261134 734 262070 856
rect 262238 734 263174 856
rect 263342 734 264278 856
rect 264446 734 265382 856
rect 265550 734 266486 856
rect 266654 734 267590 856
rect 267758 734 268694 856
rect 268862 734 269798 856
rect 269966 734 270902 856
rect 271070 734 272006 856
rect 272174 734 273110 856
rect 273278 734 274214 856
rect 274382 734 275318 856
rect 275486 734 276422 856
rect 276590 734 277526 856
rect 277694 734 278630 856
rect 278798 734 279734 856
rect 279902 734 280838 856
rect 281006 734 281942 856
rect 282110 734 283046 856
rect 283214 734 284150 856
rect 284318 734 285254 856
rect 285422 734 286358 856
rect 286526 734 287462 856
rect 287630 734 288566 856
rect 288734 734 289670 856
rect 289838 734 290774 856
rect 290942 734 291878 856
rect 292046 734 292982 856
rect 293150 734 294086 856
rect 294254 734 295190 856
rect 295358 734 296294 856
rect 296462 734 297398 856
rect 297566 734 298502 856
rect 298670 734 299606 856
rect 299774 734 300710 856
rect 300878 734 301814 856
rect 301982 734 302918 856
rect 303086 734 304022 856
rect 304190 734 305126 856
rect 305294 734 306230 856
rect 306398 734 307334 856
rect 307502 734 308438 856
rect 308606 734 309542 856
rect 309710 734 310646 856
rect 310814 734 311750 856
rect 311918 734 312854 856
rect 313022 734 313958 856
rect 314126 734 315062 856
rect 315230 734 316166 856
rect 316334 734 317270 856
rect 317438 734 318374 856
rect 318542 734 319478 856
rect 319646 734 320582 856
rect 320750 734 321686 856
rect 321854 734 322790 856
rect 322958 734 323894 856
rect 324062 734 324998 856
rect 325166 734 326102 856
rect 326270 734 327206 856
rect 327374 734 328310 856
rect 328478 734 329414 856
rect 329582 734 330518 856
rect 330686 734 331622 856
rect 331790 734 332726 856
rect 332894 734 333830 856
rect 333998 734 334934 856
rect 335102 734 336038 856
rect 336206 734 337142 856
rect 337310 734 338246 856
rect 338414 734 339350 856
rect 339518 734 340454 856
rect 340622 734 341558 856
rect 341726 734 342662 856
rect 342830 734 343766 856
rect 343934 734 344870 856
rect 345038 734 345974 856
rect 346142 734 347078 856
rect 347246 734 348182 856
rect 348350 734 349286 856
rect 349454 734 350390 856
rect 350558 734 351494 856
rect 351662 734 352598 856
rect 352766 734 353702 856
rect 353870 734 354806 856
rect 354974 734 355910 856
rect 356078 734 357014 856
rect 357182 734 358118 856
rect 358286 734 359222 856
rect 359390 734 360326 856
rect 360494 734 361430 856
rect 361598 734 362534 856
rect 362702 734 363638 856
rect 363806 734 364742 856
rect 364910 734 365846 856
rect 366014 734 366950 856
rect 367118 734 368054 856
rect 368222 734 369158 856
rect 369326 734 370262 856
rect 370430 734 371366 856
rect 371534 734 372470 856
rect 372638 734 373574 856
rect 373742 734 374678 856
rect 374846 734 375782 856
rect 375950 734 376886 856
rect 377054 734 377990 856
rect 378158 734 379094 856
rect 379262 734 380198 856
rect 380366 734 381302 856
rect 381470 734 382406 856
rect 382574 734 383510 856
rect 383678 734 384614 856
rect 384782 734 385718 856
rect 385886 734 386822 856
rect 386990 734 387926 856
rect 388094 734 389030 856
rect 389198 734 390134 856
rect 390302 734 391238 856
rect 391406 734 392342 856
rect 392510 734 393446 856
rect 393614 734 394550 856
rect 394718 734 395654 856
rect 395822 734 396758 856
rect 396926 734 397862 856
rect 398030 734 398966 856
rect 399134 734 400070 856
rect 400238 734 401174 856
rect 401342 734 402278 856
rect 402446 734 403382 856
rect 403550 734 404486 856
rect 404654 734 405590 856
rect 405758 734 406694 856
rect 406862 734 407798 856
rect 407966 734 408902 856
rect 409070 734 410006 856
rect 410174 734 411110 856
rect 411278 734 412214 856
rect 412382 734 413318 856
rect 413486 734 414422 856
rect 414590 734 415526 856
rect 415694 734 416630 856
rect 416798 734 417734 856
rect 417902 734 418838 856
rect 419006 734 419942 856
rect 420110 734 421046 856
rect 421214 734 422150 856
rect 422318 734 423254 856
rect 423422 734 424358 856
rect 424526 734 425462 856
rect 425630 734 426566 856
rect 426734 734 427670 856
rect 427838 734 428774 856
rect 428942 734 429878 856
rect 430046 734 430982 856
rect 431150 734 432086 856
rect 432254 734 433190 856
rect 433358 734 434294 856
rect 434462 734 435398 856
rect 435566 734 436502 856
rect 436670 734 437606 856
rect 437774 734 438710 856
rect 438878 734 439814 856
rect 439982 734 440918 856
rect 441086 734 442022 856
rect 442190 734 443126 856
rect 443294 734 444230 856
rect 444398 734 445334 856
rect 445502 734 446438 856
rect 446606 734 447542 856
rect 447710 734 448646 856
rect 448814 734 449750 856
rect 449918 734 450854 856
rect 451022 734 451958 856
rect 452126 734 453062 856
rect 453230 734 454166 856
rect 454334 734 455270 856
rect 455438 734 456374 856
rect 456542 734 457478 856
rect 457646 734 458582 856
rect 458750 734 459686 856
rect 459854 734 460790 856
rect 460958 734 461894 856
rect 462062 734 462998 856
rect 463166 734 464102 856
rect 464270 734 465206 856
rect 465374 734 466310 856
rect 466478 734 467414 856
rect 467582 734 468518 856
rect 468686 734 469622 856
rect 469790 734 470726 856
rect 470894 734 471830 856
rect 471998 734 472934 856
rect 473102 734 474038 856
rect 474206 734 475142 856
rect 475310 734 476246 856
rect 476414 734 477350 856
rect 477518 734 478454 856
rect 478622 734 479558 856
rect 479726 734 480662 856
rect 480830 734 481766 856
rect 481934 734 482870 856
rect 483038 734 483974 856
rect 484142 734 485078 856
rect 485246 734 486182 856
rect 486350 734 487286 856
rect 487454 734 488390 856
rect 488558 734 489494 856
rect 489662 734 490598 856
rect 490766 734 491702 856
rect 491870 734 492806 856
rect 492974 734 493910 856
rect 494078 734 495014 856
rect 495182 734 496118 856
rect 496286 734 497222 856
rect 497390 734 498326 856
rect 498494 734 499430 856
rect 499598 734 500534 856
rect 500702 734 501638 856
rect 501806 734 502742 856
rect 502910 734 503846 856
rect 504014 734 504950 856
rect 505118 734 506054 856
rect 506222 734 507158 856
rect 507326 734 508262 856
rect 508430 734 509366 856
rect 509534 734 510470 856
rect 510638 734 511574 856
rect 511742 734 512678 856
rect 512846 734 513782 856
rect 513950 734 514886 856
rect 515054 734 515990 856
rect 516158 734 517094 856
rect 517262 734 518198 856
rect 518366 734 519302 856
rect 519470 734 520406 856
rect 520574 734 521510 856
rect 521678 734 522614 856
rect 522782 734 523718 856
rect 523886 734 524822 856
rect 524990 734 525926 856
rect 526094 734 527030 856
rect 527198 734 528134 856
rect 528302 734 529238 856
rect 529406 734 530342 856
rect 530510 734 531446 856
rect 531614 734 532550 856
rect 532718 734 533654 856
rect 533822 734 534758 856
rect 534926 734 535862 856
rect 536030 734 536966 856
rect 537134 734 538070 856
rect 538238 734 539174 856
rect 539342 734 540278 856
rect 540446 734 541382 856
rect 541550 734 542486 856
rect 542654 734 543590 856
rect 543758 734 544694 856
rect 544862 734 545798 856
rect 545966 734 546902 856
rect 547070 734 548006 856
rect 548174 734 549110 856
rect 549278 734 552624 856
<< metal3 >>
rect 553404 658520 554204 658640
rect 0 657568 800 657688
rect 553404 646008 554204 646128
rect 0 645328 800 645448
rect 553404 633496 554204 633616
rect 0 633088 800 633208
rect 0 620848 800 620968
rect 553404 620984 554204 621104
rect 0 608608 800 608728
rect 553404 608472 554204 608592
rect 0 596368 800 596488
rect 553404 595960 554204 596080
rect 0 584128 800 584248
rect 553404 583448 554204 583568
rect 0 571888 800 572008
rect 553404 570936 554204 571056
rect 0 559648 800 559768
rect 553404 558424 554204 558544
rect 0 547408 800 547528
rect 553404 545912 554204 546032
rect 0 535168 800 535288
rect 553404 533400 554204 533520
rect 0 522928 800 523048
rect 553404 520888 554204 521008
rect 0 510688 800 510808
rect 553404 508376 554204 508496
rect 0 498448 800 498568
rect 553404 495864 554204 495984
rect 0 486208 800 486328
rect 553404 483352 554204 483472
rect 0 473968 800 474088
rect 553404 470840 554204 470960
rect 0 461728 800 461848
rect 553404 458328 554204 458448
rect 0 449488 800 449608
rect 553404 445816 554204 445936
rect 0 437248 800 437368
rect 553404 433304 554204 433424
rect 0 425008 800 425128
rect 553404 420792 554204 420912
rect 0 412768 800 412888
rect 553404 408280 554204 408400
rect 0 400528 800 400648
rect 553404 395768 554204 395888
rect 0 388288 800 388408
rect 553404 383256 554204 383376
rect 0 376048 800 376168
rect 553404 370744 554204 370864
rect 0 363808 800 363928
rect 553404 358232 554204 358352
rect 0 351568 800 351688
rect 553404 345720 554204 345840
rect 0 339328 800 339448
rect 553404 333208 554204 333328
rect 0 327088 800 327208
rect 553404 320696 554204 320816
rect 0 314848 800 314968
rect 553404 308184 554204 308304
rect 0 302608 800 302728
rect 553404 295672 554204 295792
rect 0 290368 800 290488
rect 553404 283160 554204 283280
rect 0 278128 800 278248
rect 553404 270648 554204 270768
rect 0 265888 800 266008
rect 553404 258136 554204 258256
rect 0 253648 800 253768
rect 553404 245624 554204 245744
rect 0 241408 800 241528
rect 553404 233112 554204 233232
rect 0 229168 800 229288
rect 553404 220600 554204 220720
rect 0 216928 800 217048
rect 553404 208088 554204 208208
rect 0 204688 800 204808
rect 553404 195576 554204 195696
rect 0 192448 800 192568
rect 553404 183064 554204 183184
rect 0 180208 800 180328
rect 553404 170552 554204 170672
rect 0 167968 800 168088
rect 553404 158040 554204 158160
rect 0 155728 800 155848
rect 553404 145528 554204 145648
rect 0 143488 800 143608
rect 553404 133016 554204 133136
rect 0 131248 800 131368
rect 553404 120504 554204 120624
rect 0 119008 800 119128
rect 553404 107992 554204 108112
rect 0 106768 800 106888
rect 553404 95480 554204 95600
rect 0 94528 800 94648
rect 553404 82968 554204 83088
rect 0 82288 800 82408
rect 553404 70456 554204 70576
rect 0 70048 800 70168
rect 0 57808 800 57928
rect 553404 57944 554204 58064
rect 0 45568 800 45688
rect 553404 45432 554204 45552
rect 0 33328 800 33448
rect 553404 32920 554204 33040
rect 0 21088 800 21208
rect 553404 20408 554204 20528
rect 0 8848 800 8968
rect 553404 7896 554204 8016
<< obsm3 >>
rect 565 658720 553404 664257
rect 565 658440 553324 658720
rect 565 657768 553404 658440
rect 880 657488 553404 657768
rect 565 646208 553404 657488
rect 565 645928 553324 646208
rect 565 645528 553404 645928
rect 880 645248 553404 645528
rect 565 633696 553404 645248
rect 565 633416 553324 633696
rect 565 633288 553404 633416
rect 880 633008 553404 633288
rect 565 621184 553404 633008
rect 565 621048 553324 621184
rect 880 620904 553324 621048
rect 880 620768 553404 620904
rect 565 608808 553404 620768
rect 880 608672 553404 608808
rect 880 608528 553324 608672
rect 565 608392 553324 608528
rect 565 596568 553404 608392
rect 880 596288 553404 596568
rect 565 596160 553404 596288
rect 565 595880 553324 596160
rect 565 584328 553404 595880
rect 880 584048 553404 584328
rect 565 583648 553404 584048
rect 565 583368 553324 583648
rect 565 572088 553404 583368
rect 880 571808 553404 572088
rect 565 571136 553404 571808
rect 565 570856 553324 571136
rect 565 559848 553404 570856
rect 880 559568 553404 559848
rect 565 558624 553404 559568
rect 565 558344 553324 558624
rect 565 547608 553404 558344
rect 880 547328 553404 547608
rect 565 546112 553404 547328
rect 565 545832 553324 546112
rect 565 535368 553404 545832
rect 880 535088 553404 535368
rect 565 533600 553404 535088
rect 565 533320 553324 533600
rect 565 523128 553404 533320
rect 880 522848 553404 523128
rect 565 521088 553404 522848
rect 565 520808 553324 521088
rect 565 510888 553404 520808
rect 880 510608 553404 510888
rect 565 508576 553404 510608
rect 565 508296 553324 508576
rect 565 498648 553404 508296
rect 880 498368 553404 498648
rect 565 496064 553404 498368
rect 565 495784 553324 496064
rect 565 486408 553404 495784
rect 880 486128 553404 486408
rect 565 483552 553404 486128
rect 565 483272 553324 483552
rect 565 474168 553404 483272
rect 880 473888 553404 474168
rect 565 471040 553404 473888
rect 565 470760 553324 471040
rect 565 461928 553404 470760
rect 880 461648 553404 461928
rect 565 458528 553404 461648
rect 565 458248 553324 458528
rect 565 449688 553404 458248
rect 880 449408 553404 449688
rect 565 446016 553404 449408
rect 565 445736 553324 446016
rect 565 437448 553404 445736
rect 880 437168 553404 437448
rect 565 433504 553404 437168
rect 565 433224 553324 433504
rect 565 425208 553404 433224
rect 880 424928 553404 425208
rect 565 420992 553404 424928
rect 565 420712 553324 420992
rect 565 412968 553404 420712
rect 880 412688 553404 412968
rect 565 408480 553404 412688
rect 565 408200 553324 408480
rect 565 400728 553404 408200
rect 880 400448 553404 400728
rect 565 395968 553404 400448
rect 565 395688 553324 395968
rect 565 388488 553404 395688
rect 880 388208 553404 388488
rect 565 383456 553404 388208
rect 565 383176 553324 383456
rect 565 376248 553404 383176
rect 880 375968 553404 376248
rect 565 370944 553404 375968
rect 565 370664 553324 370944
rect 565 364008 553404 370664
rect 880 363728 553404 364008
rect 565 358432 553404 363728
rect 565 358152 553324 358432
rect 565 351768 553404 358152
rect 880 351488 553404 351768
rect 565 345920 553404 351488
rect 565 345640 553324 345920
rect 565 339528 553404 345640
rect 880 339248 553404 339528
rect 565 333408 553404 339248
rect 565 333128 553324 333408
rect 565 327288 553404 333128
rect 880 327008 553404 327288
rect 565 320896 553404 327008
rect 565 320616 553324 320896
rect 565 315048 553404 320616
rect 880 314768 553404 315048
rect 565 308384 553404 314768
rect 565 308104 553324 308384
rect 565 302808 553404 308104
rect 880 302528 553404 302808
rect 565 295872 553404 302528
rect 565 295592 553324 295872
rect 565 290568 553404 295592
rect 880 290288 553404 290568
rect 565 283360 553404 290288
rect 565 283080 553324 283360
rect 565 278328 553404 283080
rect 880 278048 553404 278328
rect 565 270848 553404 278048
rect 565 270568 553324 270848
rect 565 266088 553404 270568
rect 880 265808 553404 266088
rect 565 258336 553404 265808
rect 565 258056 553324 258336
rect 565 253848 553404 258056
rect 880 253568 553404 253848
rect 565 245824 553404 253568
rect 565 245544 553324 245824
rect 565 241608 553404 245544
rect 880 241328 553404 241608
rect 565 233312 553404 241328
rect 565 233032 553324 233312
rect 565 229368 553404 233032
rect 880 229088 553404 229368
rect 565 220800 553404 229088
rect 565 220520 553324 220800
rect 565 217128 553404 220520
rect 880 216848 553404 217128
rect 565 208288 553404 216848
rect 565 208008 553324 208288
rect 565 204888 553404 208008
rect 880 204608 553404 204888
rect 565 195776 553404 204608
rect 565 195496 553324 195776
rect 565 192648 553404 195496
rect 880 192368 553404 192648
rect 565 183264 553404 192368
rect 565 182984 553324 183264
rect 565 180408 553404 182984
rect 880 180128 553404 180408
rect 565 170752 553404 180128
rect 565 170472 553324 170752
rect 565 168168 553404 170472
rect 880 167888 553404 168168
rect 565 158240 553404 167888
rect 565 157960 553324 158240
rect 565 155928 553404 157960
rect 880 155648 553404 155928
rect 565 145728 553404 155648
rect 565 145448 553324 145728
rect 565 143688 553404 145448
rect 880 143408 553404 143688
rect 565 133216 553404 143408
rect 565 132936 553324 133216
rect 565 131448 553404 132936
rect 880 131168 553404 131448
rect 565 120704 553404 131168
rect 565 120424 553324 120704
rect 565 119208 553404 120424
rect 880 118928 553404 119208
rect 565 108192 553404 118928
rect 565 107912 553324 108192
rect 565 106968 553404 107912
rect 880 106688 553404 106968
rect 565 95680 553404 106688
rect 565 95400 553324 95680
rect 565 94728 553404 95400
rect 880 94448 553404 94728
rect 565 83168 553404 94448
rect 565 82888 553324 83168
rect 565 82488 553404 82888
rect 880 82208 553404 82488
rect 565 70656 553404 82208
rect 565 70376 553324 70656
rect 565 70248 553404 70376
rect 880 69968 553404 70248
rect 565 58144 553404 69968
rect 565 58008 553324 58144
rect 880 57864 553324 58008
rect 880 57728 553404 57864
rect 565 45768 553404 57728
rect 880 45632 553404 45768
rect 880 45488 553324 45632
rect 565 45352 553324 45488
rect 565 33528 553404 45352
rect 880 33248 553404 33528
rect 565 33120 553404 33248
rect 565 32840 553324 33120
rect 565 21288 553404 32840
rect 880 21008 553404 21288
rect 565 20608 553404 21008
rect 565 20328 553324 20608
rect 565 9048 553404 20328
rect 880 8768 553404 9048
rect 565 8096 553404 8768
rect 565 7816 553324 8096
rect 565 2143 553404 7816
<< metal4 >>
rect 4208 2128 4528 664272
rect 19568 2128 19888 664272
rect 34928 2128 35248 664272
rect 50288 2128 50608 664272
rect 65648 2128 65968 664272
rect 81008 2128 81328 664272
rect 96368 2128 96688 664272
rect 111728 2128 112048 664272
rect 127088 2128 127408 664272
rect 142448 2128 142768 664272
rect 157808 2128 158128 664272
rect 173168 2128 173488 664272
rect 188528 2128 188848 664272
rect 203888 2128 204208 664272
rect 219248 2128 219568 664272
rect 234608 2128 234928 664272
rect 249968 2128 250288 664272
rect 265328 2128 265648 664272
rect 280688 2128 281008 664272
rect 296048 2128 296368 664272
rect 311408 2128 311728 664272
rect 326768 2128 327088 664272
rect 342128 2128 342448 664272
rect 357488 2128 357808 664272
rect 372848 2128 373168 664272
rect 388208 2128 388528 664272
rect 403568 2128 403888 664272
rect 418928 2128 419248 664272
rect 434288 2128 434608 664272
rect 449648 2128 449968 664272
rect 465008 2128 465328 664272
rect 480368 2128 480688 664272
rect 495728 2128 496048 664272
rect 511088 2128 511408 664272
rect 526448 2128 526768 664272
rect 541808 2128 542128 664272
<< obsm4 >>
rect 611 2619 4128 663917
rect 4608 2619 19488 663917
rect 19968 2619 34848 663917
rect 35328 2619 50208 663917
rect 50688 2619 65568 663917
rect 66048 2619 80928 663917
rect 81408 2619 96288 663917
rect 96768 2619 111648 663917
rect 112128 2619 127008 663917
rect 127488 2619 142368 663917
rect 142848 2619 157728 663917
rect 158208 2619 173088 663917
rect 173568 2619 188448 663917
rect 188928 2619 203808 663917
rect 204288 2619 219168 663917
rect 219648 2619 234528 663917
rect 235008 2619 249888 663917
rect 250368 2619 265248 663917
rect 265728 2619 280608 663917
rect 281088 2619 295968 663917
rect 296448 2619 311328 663917
rect 311808 2619 326688 663917
rect 327168 2619 342048 663917
rect 342528 2619 357408 663917
rect 357888 2619 372768 663917
rect 373248 2619 388128 663917
rect 388608 2619 403488 663917
rect 403968 2619 418848 663917
rect 419328 2619 434208 663917
rect 434688 2619 449568 663917
rect 450048 2619 464928 663917
rect 465408 2619 480288 663917
rect 480768 2619 495648 663917
rect 496128 2619 511008 663917
rect 511488 2619 526368 663917
rect 526848 2619 541728 663917
rect 542208 2619 551757 663917
<< labels >>
rlabel metal3 s 553404 270648 554204 270768 6 analog_io[0]
port 1 nsew signal bidirectional
rlabel metal2 s 423034 665948 423090 666748 6 analog_io[10]
port 2 nsew signal bidirectional
rlabel metal2 s 361578 665948 361634 666748 6 analog_io[11]
port 3 nsew signal bidirectional
rlabel metal2 s 300122 665948 300178 666748 6 analog_io[12]
port 4 nsew signal bidirectional
rlabel metal2 s 238666 665948 238722 666748 6 analog_io[13]
port 5 nsew signal bidirectional
rlabel metal2 s 177210 665948 177266 666748 6 analog_io[14]
port 6 nsew signal bidirectional
rlabel metal2 s 115754 665948 115810 666748 6 analog_io[15]
port 7 nsew signal bidirectional
rlabel metal2 s 54298 665948 54354 666748 6 analog_io[16]
port 8 nsew signal bidirectional
rlabel metal3 s 0 657568 800 657688 6 analog_io[17]
port 9 nsew signal bidirectional
rlabel metal3 s 0 608608 800 608728 6 analog_io[18]
port 10 nsew signal bidirectional
rlabel metal3 s 0 559648 800 559768 6 analog_io[19]
port 11 nsew signal bidirectional
rlabel metal3 s 553404 320696 554204 320816 6 analog_io[1]
port 12 nsew signal bidirectional
rlabel metal3 s 0 510688 800 510808 6 analog_io[20]
port 13 nsew signal bidirectional
rlabel metal3 s 0 461728 800 461848 6 analog_io[21]
port 14 nsew signal bidirectional
rlabel metal3 s 0 412768 800 412888 6 analog_io[22]
port 15 nsew signal bidirectional
rlabel metal3 s 0 363808 800 363928 6 analog_io[23]
port 16 nsew signal bidirectional
rlabel metal3 s 0 314848 800 314968 6 analog_io[24]
port 17 nsew signal bidirectional
rlabel metal3 s 0 265888 800 266008 6 analog_io[25]
port 18 nsew signal bidirectional
rlabel metal3 s 0 216928 800 217048 6 analog_io[26]
port 19 nsew signal bidirectional
rlabel metal3 s 0 167968 800 168088 6 analog_io[27]
port 20 nsew signal bidirectional
rlabel metal3 s 0 119008 800 119128 6 analog_io[28]
port 21 nsew signal bidirectional
rlabel metal3 s 553404 370744 554204 370864 6 analog_io[2]
port 22 nsew signal bidirectional
rlabel metal3 s 553404 420792 554204 420912 6 analog_io[3]
port 23 nsew signal bidirectional
rlabel metal3 s 553404 470840 554204 470960 6 analog_io[4]
port 24 nsew signal bidirectional
rlabel metal3 s 553404 520888 554204 521008 6 analog_io[5]
port 25 nsew signal bidirectional
rlabel metal3 s 553404 570936 554204 571056 6 analog_io[6]
port 26 nsew signal bidirectional
rlabel metal3 s 553404 620984 554204 621104 6 analog_io[7]
port 27 nsew signal bidirectional
rlabel metal2 s 545946 665948 546002 666748 6 analog_io[8]
port 28 nsew signal bidirectional
rlabel metal2 s 484490 665948 484546 666748 6 analog_io[9]
port 29 nsew signal bidirectional
rlabel metal3 s 553404 7896 554204 8016 6 io_in[0]
port 30 nsew signal input
rlabel metal3 s 553404 433304 554204 433424 6 io_in[10]
port 31 nsew signal input
rlabel metal3 s 553404 483352 554204 483472 6 io_in[11]
port 32 nsew signal input
rlabel metal3 s 553404 533400 554204 533520 6 io_in[12]
port 33 nsew signal input
rlabel metal3 s 553404 583448 554204 583568 6 io_in[13]
port 34 nsew signal input
rlabel metal3 s 553404 633496 554204 633616 6 io_in[14]
port 35 nsew signal input
rlabel metal2 s 530582 665948 530638 666748 6 io_in[15]
port 36 nsew signal input
rlabel metal2 s 469126 665948 469182 666748 6 io_in[16]
port 37 nsew signal input
rlabel metal2 s 407670 665948 407726 666748 6 io_in[17]
port 38 nsew signal input
rlabel metal2 s 346214 665948 346270 666748 6 io_in[18]
port 39 nsew signal input
rlabel metal2 s 284758 665948 284814 666748 6 io_in[19]
port 40 nsew signal input
rlabel metal3 s 553404 45432 554204 45552 6 io_in[1]
port 41 nsew signal input
rlabel metal2 s 223302 665948 223358 666748 6 io_in[20]
port 42 nsew signal input
rlabel metal2 s 161846 665948 161902 666748 6 io_in[21]
port 43 nsew signal input
rlabel metal2 s 100390 665948 100446 666748 6 io_in[22]
port 44 nsew signal input
rlabel metal2 s 38934 665948 38990 666748 6 io_in[23]
port 45 nsew signal input
rlabel metal3 s 0 645328 800 645448 6 io_in[24]
port 46 nsew signal input
rlabel metal3 s 0 596368 800 596488 6 io_in[25]
port 47 nsew signal input
rlabel metal3 s 0 547408 800 547528 6 io_in[26]
port 48 nsew signal input
rlabel metal3 s 0 498448 800 498568 6 io_in[27]
port 49 nsew signal input
rlabel metal3 s 0 449488 800 449608 6 io_in[28]
port 50 nsew signal input
rlabel metal3 s 0 400528 800 400648 6 io_in[29]
port 51 nsew signal input
rlabel metal3 s 553404 82968 554204 83088 6 io_in[2]
port 52 nsew signal input
rlabel metal3 s 0 351568 800 351688 6 io_in[30]
port 53 nsew signal input
rlabel metal3 s 0 302608 800 302728 6 io_in[31]
port 54 nsew signal input
rlabel metal3 s 0 253648 800 253768 6 io_in[32]
port 55 nsew signal input
rlabel metal3 s 0 204688 800 204808 6 io_in[33]
port 56 nsew signal input
rlabel metal3 s 0 155728 800 155848 6 io_in[34]
port 57 nsew signal input
rlabel metal3 s 0 106768 800 106888 6 io_in[35]
port 58 nsew signal input
rlabel metal3 s 0 70048 800 70168 6 io_in[36]
port 59 nsew signal input
rlabel metal3 s 0 33328 800 33448 6 io_in[37]
port 60 nsew signal input
rlabel metal3 s 553404 120504 554204 120624 6 io_in[3]
port 61 nsew signal input
rlabel metal3 s 553404 158040 554204 158160 6 io_in[4]
port 62 nsew signal input
rlabel metal3 s 553404 195576 554204 195696 6 io_in[5]
port 63 nsew signal input
rlabel metal3 s 553404 233112 554204 233232 6 io_in[6]
port 64 nsew signal input
rlabel metal3 s 553404 283160 554204 283280 6 io_in[7]
port 65 nsew signal input
rlabel metal3 s 553404 333208 554204 333328 6 io_in[8]
port 66 nsew signal input
rlabel metal3 s 553404 383256 554204 383376 6 io_in[9]
port 67 nsew signal input
rlabel metal3 s 553404 32920 554204 33040 6 io_oeb[0]
port 68 nsew signal output
rlabel metal3 s 553404 458328 554204 458448 6 io_oeb[10]
port 69 nsew signal output
rlabel metal3 s 553404 508376 554204 508496 6 io_oeb[11]
port 70 nsew signal output
rlabel metal3 s 553404 558424 554204 558544 6 io_oeb[12]
port 71 nsew signal output
rlabel metal3 s 553404 608472 554204 608592 6 io_oeb[13]
port 72 nsew signal output
rlabel metal3 s 553404 658520 554204 658640 6 io_oeb[14]
port 73 nsew signal output
rlabel metal2 s 499854 665948 499910 666748 6 io_oeb[15]
port 74 nsew signal output
rlabel metal2 s 438398 665948 438454 666748 6 io_oeb[16]
port 75 nsew signal output
rlabel metal2 s 376942 665948 376998 666748 6 io_oeb[17]
port 76 nsew signal output
rlabel metal2 s 315486 665948 315542 666748 6 io_oeb[18]
port 77 nsew signal output
rlabel metal2 s 254030 665948 254086 666748 6 io_oeb[19]
port 78 nsew signal output
rlabel metal3 s 553404 70456 554204 70576 6 io_oeb[1]
port 79 nsew signal output
rlabel metal2 s 192574 665948 192630 666748 6 io_oeb[20]
port 80 nsew signal output
rlabel metal2 s 131118 665948 131174 666748 6 io_oeb[21]
port 81 nsew signal output
rlabel metal2 s 69662 665948 69718 666748 6 io_oeb[22]
port 82 nsew signal output
rlabel metal2 s 8206 665948 8262 666748 6 io_oeb[23]
port 83 nsew signal output
rlabel metal3 s 0 620848 800 620968 6 io_oeb[24]
port 84 nsew signal output
rlabel metal3 s 0 571888 800 572008 6 io_oeb[25]
port 85 nsew signal output
rlabel metal3 s 0 522928 800 523048 6 io_oeb[26]
port 86 nsew signal output
rlabel metal3 s 0 473968 800 474088 6 io_oeb[27]
port 87 nsew signal output
rlabel metal3 s 0 425008 800 425128 6 io_oeb[28]
port 88 nsew signal output
rlabel metal3 s 0 376048 800 376168 6 io_oeb[29]
port 89 nsew signal output
rlabel metal3 s 553404 107992 554204 108112 6 io_oeb[2]
port 90 nsew signal output
rlabel metal3 s 0 327088 800 327208 6 io_oeb[30]
port 91 nsew signal output
rlabel metal3 s 0 278128 800 278248 6 io_oeb[31]
port 92 nsew signal output
rlabel metal3 s 0 229168 800 229288 6 io_oeb[32]
port 93 nsew signal output
rlabel metal3 s 0 180208 800 180328 6 io_oeb[33]
port 94 nsew signal output
rlabel metal3 s 0 131248 800 131368 6 io_oeb[34]
port 95 nsew signal output
rlabel metal3 s 0 82288 800 82408 6 io_oeb[35]
port 96 nsew signal output
rlabel metal3 s 0 45568 800 45688 6 io_oeb[36]
port 97 nsew signal output
rlabel metal3 s 0 8848 800 8968 6 io_oeb[37]
port 98 nsew signal output
rlabel metal3 s 553404 145528 554204 145648 6 io_oeb[3]
port 99 nsew signal output
rlabel metal3 s 553404 183064 554204 183184 6 io_oeb[4]
port 100 nsew signal output
rlabel metal3 s 553404 220600 554204 220720 6 io_oeb[5]
port 101 nsew signal output
rlabel metal3 s 553404 258136 554204 258256 6 io_oeb[6]
port 102 nsew signal output
rlabel metal3 s 553404 308184 554204 308304 6 io_oeb[7]
port 103 nsew signal output
rlabel metal3 s 553404 358232 554204 358352 6 io_oeb[8]
port 104 nsew signal output
rlabel metal3 s 553404 408280 554204 408400 6 io_oeb[9]
port 105 nsew signal output
rlabel metal3 s 553404 20408 554204 20528 6 io_out[0]
port 106 nsew signal output
rlabel metal3 s 553404 445816 554204 445936 6 io_out[10]
port 107 nsew signal output
rlabel metal3 s 553404 495864 554204 495984 6 io_out[11]
port 108 nsew signal output
rlabel metal3 s 553404 545912 554204 546032 6 io_out[12]
port 109 nsew signal output
rlabel metal3 s 553404 595960 554204 596080 6 io_out[13]
port 110 nsew signal output
rlabel metal3 s 553404 646008 554204 646128 6 io_out[14]
port 111 nsew signal output
rlabel metal2 s 515218 665948 515274 666748 6 io_out[15]
port 112 nsew signal output
rlabel metal2 s 453762 665948 453818 666748 6 io_out[16]
port 113 nsew signal output
rlabel metal2 s 392306 665948 392362 666748 6 io_out[17]
port 114 nsew signal output
rlabel metal2 s 330850 665948 330906 666748 6 io_out[18]
port 115 nsew signal output
rlabel metal2 s 269394 665948 269450 666748 6 io_out[19]
port 116 nsew signal output
rlabel metal3 s 553404 57944 554204 58064 6 io_out[1]
port 117 nsew signal output
rlabel metal2 s 207938 665948 207994 666748 6 io_out[20]
port 118 nsew signal output
rlabel metal2 s 146482 665948 146538 666748 6 io_out[21]
port 119 nsew signal output
rlabel metal2 s 85026 665948 85082 666748 6 io_out[22]
port 120 nsew signal output
rlabel metal2 s 23570 665948 23626 666748 6 io_out[23]
port 121 nsew signal output
rlabel metal3 s 0 633088 800 633208 6 io_out[24]
port 122 nsew signal output
rlabel metal3 s 0 584128 800 584248 6 io_out[25]
port 123 nsew signal output
rlabel metal3 s 0 535168 800 535288 6 io_out[26]
port 124 nsew signal output
rlabel metal3 s 0 486208 800 486328 6 io_out[27]
port 125 nsew signal output
rlabel metal3 s 0 437248 800 437368 6 io_out[28]
port 126 nsew signal output
rlabel metal3 s 0 388288 800 388408 6 io_out[29]
port 127 nsew signal output
rlabel metal3 s 553404 95480 554204 95600 6 io_out[2]
port 128 nsew signal output
rlabel metal3 s 0 339328 800 339448 6 io_out[30]
port 129 nsew signal output
rlabel metal3 s 0 290368 800 290488 6 io_out[31]
port 130 nsew signal output
rlabel metal3 s 0 241408 800 241528 6 io_out[32]
port 131 nsew signal output
rlabel metal3 s 0 192448 800 192568 6 io_out[33]
port 132 nsew signal output
rlabel metal3 s 0 143488 800 143608 6 io_out[34]
port 133 nsew signal output
rlabel metal3 s 0 94528 800 94648 6 io_out[35]
port 134 nsew signal output
rlabel metal3 s 0 57808 800 57928 6 io_out[36]
port 135 nsew signal output
rlabel metal3 s 0 21088 800 21208 6 io_out[37]
port 136 nsew signal output
rlabel metal3 s 553404 133016 554204 133136 6 io_out[3]
port 137 nsew signal output
rlabel metal3 s 553404 170552 554204 170672 6 io_out[4]
port 138 nsew signal output
rlabel metal3 s 553404 208088 554204 208208 6 io_out[5]
port 139 nsew signal output
rlabel metal3 s 553404 245624 554204 245744 6 io_out[6]
port 140 nsew signal output
rlabel metal3 s 553404 295672 554204 295792 6 io_out[7]
port 141 nsew signal output
rlabel metal3 s 553404 345720 554204 345840 6 io_out[8]
port 142 nsew signal output
rlabel metal3 s 553404 395768 554204 395888 6 io_out[9]
port 143 nsew signal output
rlabel metal2 s 121918 0 121974 800 6 la_data_in[0]
port 144 nsew signal input
rlabel metal2 s 453118 0 453174 800 6 la_data_in[100]
port 145 nsew signal input
rlabel metal2 s 456430 0 456486 800 6 la_data_in[101]
port 146 nsew signal input
rlabel metal2 s 459742 0 459798 800 6 la_data_in[102]
port 147 nsew signal input
rlabel metal2 s 463054 0 463110 800 6 la_data_in[103]
port 148 nsew signal input
rlabel metal2 s 466366 0 466422 800 6 la_data_in[104]
port 149 nsew signal input
rlabel metal2 s 469678 0 469734 800 6 la_data_in[105]
port 150 nsew signal input
rlabel metal2 s 472990 0 473046 800 6 la_data_in[106]
port 151 nsew signal input
rlabel metal2 s 476302 0 476358 800 6 la_data_in[107]
port 152 nsew signal input
rlabel metal2 s 479614 0 479670 800 6 la_data_in[108]
port 153 nsew signal input
rlabel metal2 s 482926 0 482982 800 6 la_data_in[109]
port 154 nsew signal input
rlabel metal2 s 155038 0 155094 800 6 la_data_in[10]
port 155 nsew signal input
rlabel metal2 s 486238 0 486294 800 6 la_data_in[110]
port 156 nsew signal input
rlabel metal2 s 489550 0 489606 800 6 la_data_in[111]
port 157 nsew signal input
rlabel metal2 s 492862 0 492918 800 6 la_data_in[112]
port 158 nsew signal input
rlabel metal2 s 496174 0 496230 800 6 la_data_in[113]
port 159 nsew signal input
rlabel metal2 s 499486 0 499542 800 6 la_data_in[114]
port 160 nsew signal input
rlabel metal2 s 502798 0 502854 800 6 la_data_in[115]
port 161 nsew signal input
rlabel metal2 s 506110 0 506166 800 6 la_data_in[116]
port 162 nsew signal input
rlabel metal2 s 509422 0 509478 800 6 la_data_in[117]
port 163 nsew signal input
rlabel metal2 s 512734 0 512790 800 6 la_data_in[118]
port 164 nsew signal input
rlabel metal2 s 516046 0 516102 800 6 la_data_in[119]
port 165 nsew signal input
rlabel metal2 s 158350 0 158406 800 6 la_data_in[11]
port 166 nsew signal input
rlabel metal2 s 519358 0 519414 800 6 la_data_in[120]
port 167 nsew signal input
rlabel metal2 s 522670 0 522726 800 6 la_data_in[121]
port 168 nsew signal input
rlabel metal2 s 525982 0 526038 800 6 la_data_in[122]
port 169 nsew signal input
rlabel metal2 s 529294 0 529350 800 6 la_data_in[123]
port 170 nsew signal input
rlabel metal2 s 532606 0 532662 800 6 la_data_in[124]
port 171 nsew signal input
rlabel metal2 s 535918 0 535974 800 6 la_data_in[125]
port 172 nsew signal input
rlabel metal2 s 539230 0 539286 800 6 la_data_in[126]
port 173 nsew signal input
rlabel metal2 s 542542 0 542598 800 6 la_data_in[127]
port 174 nsew signal input
rlabel metal2 s 161662 0 161718 800 6 la_data_in[12]
port 175 nsew signal input
rlabel metal2 s 164974 0 165030 800 6 la_data_in[13]
port 176 nsew signal input
rlabel metal2 s 168286 0 168342 800 6 la_data_in[14]
port 177 nsew signal input
rlabel metal2 s 171598 0 171654 800 6 la_data_in[15]
port 178 nsew signal input
rlabel metal2 s 174910 0 174966 800 6 la_data_in[16]
port 179 nsew signal input
rlabel metal2 s 178222 0 178278 800 6 la_data_in[17]
port 180 nsew signal input
rlabel metal2 s 181534 0 181590 800 6 la_data_in[18]
port 181 nsew signal input
rlabel metal2 s 184846 0 184902 800 6 la_data_in[19]
port 182 nsew signal input
rlabel metal2 s 125230 0 125286 800 6 la_data_in[1]
port 183 nsew signal input
rlabel metal2 s 188158 0 188214 800 6 la_data_in[20]
port 184 nsew signal input
rlabel metal2 s 191470 0 191526 800 6 la_data_in[21]
port 185 nsew signal input
rlabel metal2 s 194782 0 194838 800 6 la_data_in[22]
port 186 nsew signal input
rlabel metal2 s 198094 0 198150 800 6 la_data_in[23]
port 187 nsew signal input
rlabel metal2 s 201406 0 201462 800 6 la_data_in[24]
port 188 nsew signal input
rlabel metal2 s 204718 0 204774 800 6 la_data_in[25]
port 189 nsew signal input
rlabel metal2 s 208030 0 208086 800 6 la_data_in[26]
port 190 nsew signal input
rlabel metal2 s 211342 0 211398 800 6 la_data_in[27]
port 191 nsew signal input
rlabel metal2 s 214654 0 214710 800 6 la_data_in[28]
port 192 nsew signal input
rlabel metal2 s 217966 0 218022 800 6 la_data_in[29]
port 193 nsew signal input
rlabel metal2 s 128542 0 128598 800 6 la_data_in[2]
port 194 nsew signal input
rlabel metal2 s 221278 0 221334 800 6 la_data_in[30]
port 195 nsew signal input
rlabel metal2 s 224590 0 224646 800 6 la_data_in[31]
port 196 nsew signal input
rlabel metal2 s 227902 0 227958 800 6 la_data_in[32]
port 197 nsew signal input
rlabel metal2 s 231214 0 231270 800 6 la_data_in[33]
port 198 nsew signal input
rlabel metal2 s 234526 0 234582 800 6 la_data_in[34]
port 199 nsew signal input
rlabel metal2 s 237838 0 237894 800 6 la_data_in[35]
port 200 nsew signal input
rlabel metal2 s 241150 0 241206 800 6 la_data_in[36]
port 201 nsew signal input
rlabel metal2 s 244462 0 244518 800 6 la_data_in[37]
port 202 nsew signal input
rlabel metal2 s 247774 0 247830 800 6 la_data_in[38]
port 203 nsew signal input
rlabel metal2 s 251086 0 251142 800 6 la_data_in[39]
port 204 nsew signal input
rlabel metal2 s 131854 0 131910 800 6 la_data_in[3]
port 205 nsew signal input
rlabel metal2 s 254398 0 254454 800 6 la_data_in[40]
port 206 nsew signal input
rlabel metal2 s 257710 0 257766 800 6 la_data_in[41]
port 207 nsew signal input
rlabel metal2 s 261022 0 261078 800 6 la_data_in[42]
port 208 nsew signal input
rlabel metal2 s 264334 0 264390 800 6 la_data_in[43]
port 209 nsew signal input
rlabel metal2 s 267646 0 267702 800 6 la_data_in[44]
port 210 nsew signal input
rlabel metal2 s 270958 0 271014 800 6 la_data_in[45]
port 211 nsew signal input
rlabel metal2 s 274270 0 274326 800 6 la_data_in[46]
port 212 nsew signal input
rlabel metal2 s 277582 0 277638 800 6 la_data_in[47]
port 213 nsew signal input
rlabel metal2 s 280894 0 280950 800 6 la_data_in[48]
port 214 nsew signal input
rlabel metal2 s 284206 0 284262 800 6 la_data_in[49]
port 215 nsew signal input
rlabel metal2 s 135166 0 135222 800 6 la_data_in[4]
port 216 nsew signal input
rlabel metal2 s 287518 0 287574 800 6 la_data_in[50]
port 217 nsew signal input
rlabel metal2 s 290830 0 290886 800 6 la_data_in[51]
port 218 nsew signal input
rlabel metal2 s 294142 0 294198 800 6 la_data_in[52]
port 219 nsew signal input
rlabel metal2 s 297454 0 297510 800 6 la_data_in[53]
port 220 nsew signal input
rlabel metal2 s 300766 0 300822 800 6 la_data_in[54]
port 221 nsew signal input
rlabel metal2 s 304078 0 304134 800 6 la_data_in[55]
port 222 nsew signal input
rlabel metal2 s 307390 0 307446 800 6 la_data_in[56]
port 223 nsew signal input
rlabel metal2 s 310702 0 310758 800 6 la_data_in[57]
port 224 nsew signal input
rlabel metal2 s 314014 0 314070 800 6 la_data_in[58]
port 225 nsew signal input
rlabel metal2 s 317326 0 317382 800 6 la_data_in[59]
port 226 nsew signal input
rlabel metal2 s 138478 0 138534 800 6 la_data_in[5]
port 227 nsew signal input
rlabel metal2 s 320638 0 320694 800 6 la_data_in[60]
port 228 nsew signal input
rlabel metal2 s 323950 0 324006 800 6 la_data_in[61]
port 229 nsew signal input
rlabel metal2 s 327262 0 327318 800 6 la_data_in[62]
port 230 nsew signal input
rlabel metal2 s 330574 0 330630 800 6 la_data_in[63]
port 231 nsew signal input
rlabel metal2 s 333886 0 333942 800 6 la_data_in[64]
port 232 nsew signal input
rlabel metal2 s 337198 0 337254 800 6 la_data_in[65]
port 233 nsew signal input
rlabel metal2 s 340510 0 340566 800 6 la_data_in[66]
port 234 nsew signal input
rlabel metal2 s 343822 0 343878 800 6 la_data_in[67]
port 235 nsew signal input
rlabel metal2 s 347134 0 347190 800 6 la_data_in[68]
port 236 nsew signal input
rlabel metal2 s 350446 0 350502 800 6 la_data_in[69]
port 237 nsew signal input
rlabel metal2 s 141790 0 141846 800 6 la_data_in[6]
port 238 nsew signal input
rlabel metal2 s 353758 0 353814 800 6 la_data_in[70]
port 239 nsew signal input
rlabel metal2 s 357070 0 357126 800 6 la_data_in[71]
port 240 nsew signal input
rlabel metal2 s 360382 0 360438 800 6 la_data_in[72]
port 241 nsew signal input
rlabel metal2 s 363694 0 363750 800 6 la_data_in[73]
port 242 nsew signal input
rlabel metal2 s 367006 0 367062 800 6 la_data_in[74]
port 243 nsew signal input
rlabel metal2 s 370318 0 370374 800 6 la_data_in[75]
port 244 nsew signal input
rlabel metal2 s 373630 0 373686 800 6 la_data_in[76]
port 245 nsew signal input
rlabel metal2 s 376942 0 376998 800 6 la_data_in[77]
port 246 nsew signal input
rlabel metal2 s 380254 0 380310 800 6 la_data_in[78]
port 247 nsew signal input
rlabel metal2 s 383566 0 383622 800 6 la_data_in[79]
port 248 nsew signal input
rlabel metal2 s 145102 0 145158 800 6 la_data_in[7]
port 249 nsew signal input
rlabel metal2 s 386878 0 386934 800 6 la_data_in[80]
port 250 nsew signal input
rlabel metal2 s 390190 0 390246 800 6 la_data_in[81]
port 251 nsew signal input
rlabel metal2 s 393502 0 393558 800 6 la_data_in[82]
port 252 nsew signal input
rlabel metal2 s 396814 0 396870 800 6 la_data_in[83]
port 253 nsew signal input
rlabel metal2 s 400126 0 400182 800 6 la_data_in[84]
port 254 nsew signal input
rlabel metal2 s 403438 0 403494 800 6 la_data_in[85]
port 255 nsew signal input
rlabel metal2 s 406750 0 406806 800 6 la_data_in[86]
port 256 nsew signal input
rlabel metal2 s 410062 0 410118 800 6 la_data_in[87]
port 257 nsew signal input
rlabel metal2 s 413374 0 413430 800 6 la_data_in[88]
port 258 nsew signal input
rlabel metal2 s 416686 0 416742 800 6 la_data_in[89]
port 259 nsew signal input
rlabel metal2 s 148414 0 148470 800 6 la_data_in[8]
port 260 nsew signal input
rlabel metal2 s 419998 0 420054 800 6 la_data_in[90]
port 261 nsew signal input
rlabel metal2 s 423310 0 423366 800 6 la_data_in[91]
port 262 nsew signal input
rlabel metal2 s 426622 0 426678 800 6 la_data_in[92]
port 263 nsew signal input
rlabel metal2 s 429934 0 429990 800 6 la_data_in[93]
port 264 nsew signal input
rlabel metal2 s 433246 0 433302 800 6 la_data_in[94]
port 265 nsew signal input
rlabel metal2 s 436558 0 436614 800 6 la_data_in[95]
port 266 nsew signal input
rlabel metal2 s 439870 0 439926 800 6 la_data_in[96]
port 267 nsew signal input
rlabel metal2 s 443182 0 443238 800 6 la_data_in[97]
port 268 nsew signal input
rlabel metal2 s 446494 0 446550 800 6 la_data_in[98]
port 269 nsew signal input
rlabel metal2 s 449806 0 449862 800 6 la_data_in[99]
port 270 nsew signal input
rlabel metal2 s 151726 0 151782 800 6 la_data_in[9]
port 271 nsew signal input
rlabel metal2 s 123022 0 123078 800 6 la_data_out[0]
port 272 nsew signal output
rlabel metal2 s 454222 0 454278 800 6 la_data_out[100]
port 273 nsew signal output
rlabel metal2 s 457534 0 457590 800 6 la_data_out[101]
port 274 nsew signal output
rlabel metal2 s 460846 0 460902 800 6 la_data_out[102]
port 275 nsew signal output
rlabel metal2 s 464158 0 464214 800 6 la_data_out[103]
port 276 nsew signal output
rlabel metal2 s 467470 0 467526 800 6 la_data_out[104]
port 277 nsew signal output
rlabel metal2 s 470782 0 470838 800 6 la_data_out[105]
port 278 nsew signal output
rlabel metal2 s 474094 0 474150 800 6 la_data_out[106]
port 279 nsew signal output
rlabel metal2 s 477406 0 477462 800 6 la_data_out[107]
port 280 nsew signal output
rlabel metal2 s 480718 0 480774 800 6 la_data_out[108]
port 281 nsew signal output
rlabel metal2 s 484030 0 484086 800 6 la_data_out[109]
port 282 nsew signal output
rlabel metal2 s 156142 0 156198 800 6 la_data_out[10]
port 283 nsew signal output
rlabel metal2 s 487342 0 487398 800 6 la_data_out[110]
port 284 nsew signal output
rlabel metal2 s 490654 0 490710 800 6 la_data_out[111]
port 285 nsew signal output
rlabel metal2 s 493966 0 494022 800 6 la_data_out[112]
port 286 nsew signal output
rlabel metal2 s 497278 0 497334 800 6 la_data_out[113]
port 287 nsew signal output
rlabel metal2 s 500590 0 500646 800 6 la_data_out[114]
port 288 nsew signal output
rlabel metal2 s 503902 0 503958 800 6 la_data_out[115]
port 289 nsew signal output
rlabel metal2 s 507214 0 507270 800 6 la_data_out[116]
port 290 nsew signal output
rlabel metal2 s 510526 0 510582 800 6 la_data_out[117]
port 291 nsew signal output
rlabel metal2 s 513838 0 513894 800 6 la_data_out[118]
port 292 nsew signal output
rlabel metal2 s 517150 0 517206 800 6 la_data_out[119]
port 293 nsew signal output
rlabel metal2 s 159454 0 159510 800 6 la_data_out[11]
port 294 nsew signal output
rlabel metal2 s 520462 0 520518 800 6 la_data_out[120]
port 295 nsew signal output
rlabel metal2 s 523774 0 523830 800 6 la_data_out[121]
port 296 nsew signal output
rlabel metal2 s 527086 0 527142 800 6 la_data_out[122]
port 297 nsew signal output
rlabel metal2 s 530398 0 530454 800 6 la_data_out[123]
port 298 nsew signal output
rlabel metal2 s 533710 0 533766 800 6 la_data_out[124]
port 299 nsew signal output
rlabel metal2 s 537022 0 537078 800 6 la_data_out[125]
port 300 nsew signal output
rlabel metal2 s 540334 0 540390 800 6 la_data_out[126]
port 301 nsew signal output
rlabel metal2 s 543646 0 543702 800 6 la_data_out[127]
port 302 nsew signal output
rlabel metal2 s 162766 0 162822 800 6 la_data_out[12]
port 303 nsew signal output
rlabel metal2 s 166078 0 166134 800 6 la_data_out[13]
port 304 nsew signal output
rlabel metal2 s 169390 0 169446 800 6 la_data_out[14]
port 305 nsew signal output
rlabel metal2 s 172702 0 172758 800 6 la_data_out[15]
port 306 nsew signal output
rlabel metal2 s 176014 0 176070 800 6 la_data_out[16]
port 307 nsew signal output
rlabel metal2 s 179326 0 179382 800 6 la_data_out[17]
port 308 nsew signal output
rlabel metal2 s 182638 0 182694 800 6 la_data_out[18]
port 309 nsew signal output
rlabel metal2 s 185950 0 186006 800 6 la_data_out[19]
port 310 nsew signal output
rlabel metal2 s 126334 0 126390 800 6 la_data_out[1]
port 311 nsew signal output
rlabel metal2 s 189262 0 189318 800 6 la_data_out[20]
port 312 nsew signal output
rlabel metal2 s 192574 0 192630 800 6 la_data_out[21]
port 313 nsew signal output
rlabel metal2 s 195886 0 195942 800 6 la_data_out[22]
port 314 nsew signal output
rlabel metal2 s 199198 0 199254 800 6 la_data_out[23]
port 315 nsew signal output
rlabel metal2 s 202510 0 202566 800 6 la_data_out[24]
port 316 nsew signal output
rlabel metal2 s 205822 0 205878 800 6 la_data_out[25]
port 317 nsew signal output
rlabel metal2 s 209134 0 209190 800 6 la_data_out[26]
port 318 nsew signal output
rlabel metal2 s 212446 0 212502 800 6 la_data_out[27]
port 319 nsew signal output
rlabel metal2 s 215758 0 215814 800 6 la_data_out[28]
port 320 nsew signal output
rlabel metal2 s 219070 0 219126 800 6 la_data_out[29]
port 321 nsew signal output
rlabel metal2 s 129646 0 129702 800 6 la_data_out[2]
port 322 nsew signal output
rlabel metal2 s 222382 0 222438 800 6 la_data_out[30]
port 323 nsew signal output
rlabel metal2 s 225694 0 225750 800 6 la_data_out[31]
port 324 nsew signal output
rlabel metal2 s 229006 0 229062 800 6 la_data_out[32]
port 325 nsew signal output
rlabel metal2 s 232318 0 232374 800 6 la_data_out[33]
port 326 nsew signal output
rlabel metal2 s 235630 0 235686 800 6 la_data_out[34]
port 327 nsew signal output
rlabel metal2 s 238942 0 238998 800 6 la_data_out[35]
port 328 nsew signal output
rlabel metal2 s 242254 0 242310 800 6 la_data_out[36]
port 329 nsew signal output
rlabel metal2 s 245566 0 245622 800 6 la_data_out[37]
port 330 nsew signal output
rlabel metal2 s 248878 0 248934 800 6 la_data_out[38]
port 331 nsew signal output
rlabel metal2 s 252190 0 252246 800 6 la_data_out[39]
port 332 nsew signal output
rlabel metal2 s 132958 0 133014 800 6 la_data_out[3]
port 333 nsew signal output
rlabel metal2 s 255502 0 255558 800 6 la_data_out[40]
port 334 nsew signal output
rlabel metal2 s 258814 0 258870 800 6 la_data_out[41]
port 335 nsew signal output
rlabel metal2 s 262126 0 262182 800 6 la_data_out[42]
port 336 nsew signal output
rlabel metal2 s 265438 0 265494 800 6 la_data_out[43]
port 337 nsew signal output
rlabel metal2 s 268750 0 268806 800 6 la_data_out[44]
port 338 nsew signal output
rlabel metal2 s 272062 0 272118 800 6 la_data_out[45]
port 339 nsew signal output
rlabel metal2 s 275374 0 275430 800 6 la_data_out[46]
port 340 nsew signal output
rlabel metal2 s 278686 0 278742 800 6 la_data_out[47]
port 341 nsew signal output
rlabel metal2 s 281998 0 282054 800 6 la_data_out[48]
port 342 nsew signal output
rlabel metal2 s 285310 0 285366 800 6 la_data_out[49]
port 343 nsew signal output
rlabel metal2 s 136270 0 136326 800 6 la_data_out[4]
port 344 nsew signal output
rlabel metal2 s 288622 0 288678 800 6 la_data_out[50]
port 345 nsew signal output
rlabel metal2 s 291934 0 291990 800 6 la_data_out[51]
port 346 nsew signal output
rlabel metal2 s 295246 0 295302 800 6 la_data_out[52]
port 347 nsew signal output
rlabel metal2 s 298558 0 298614 800 6 la_data_out[53]
port 348 nsew signal output
rlabel metal2 s 301870 0 301926 800 6 la_data_out[54]
port 349 nsew signal output
rlabel metal2 s 305182 0 305238 800 6 la_data_out[55]
port 350 nsew signal output
rlabel metal2 s 308494 0 308550 800 6 la_data_out[56]
port 351 nsew signal output
rlabel metal2 s 311806 0 311862 800 6 la_data_out[57]
port 352 nsew signal output
rlabel metal2 s 315118 0 315174 800 6 la_data_out[58]
port 353 nsew signal output
rlabel metal2 s 318430 0 318486 800 6 la_data_out[59]
port 354 nsew signal output
rlabel metal2 s 139582 0 139638 800 6 la_data_out[5]
port 355 nsew signal output
rlabel metal2 s 321742 0 321798 800 6 la_data_out[60]
port 356 nsew signal output
rlabel metal2 s 325054 0 325110 800 6 la_data_out[61]
port 357 nsew signal output
rlabel metal2 s 328366 0 328422 800 6 la_data_out[62]
port 358 nsew signal output
rlabel metal2 s 331678 0 331734 800 6 la_data_out[63]
port 359 nsew signal output
rlabel metal2 s 334990 0 335046 800 6 la_data_out[64]
port 360 nsew signal output
rlabel metal2 s 338302 0 338358 800 6 la_data_out[65]
port 361 nsew signal output
rlabel metal2 s 341614 0 341670 800 6 la_data_out[66]
port 362 nsew signal output
rlabel metal2 s 344926 0 344982 800 6 la_data_out[67]
port 363 nsew signal output
rlabel metal2 s 348238 0 348294 800 6 la_data_out[68]
port 364 nsew signal output
rlabel metal2 s 351550 0 351606 800 6 la_data_out[69]
port 365 nsew signal output
rlabel metal2 s 142894 0 142950 800 6 la_data_out[6]
port 366 nsew signal output
rlabel metal2 s 354862 0 354918 800 6 la_data_out[70]
port 367 nsew signal output
rlabel metal2 s 358174 0 358230 800 6 la_data_out[71]
port 368 nsew signal output
rlabel metal2 s 361486 0 361542 800 6 la_data_out[72]
port 369 nsew signal output
rlabel metal2 s 364798 0 364854 800 6 la_data_out[73]
port 370 nsew signal output
rlabel metal2 s 368110 0 368166 800 6 la_data_out[74]
port 371 nsew signal output
rlabel metal2 s 371422 0 371478 800 6 la_data_out[75]
port 372 nsew signal output
rlabel metal2 s 374734 0 374790 800 6 la_data_out[76]
port 373 nsew signal output
rlabel metal2 s 378046 0 378102 800 6 la_data_out[77]
port 374 nsew signal output
rlabel metal2 s 381358 0 381414 800 6 la_data_out[78]
port 375 nsew signal output
rlabel metal2 s 384670 0 384726 800 6 la_data_out[79]
port 376 nsew signal output
rlabel metal2 s 146206 0 146262 800 6 la_data_out[7]
port 377 nsew signal output
rlabel metal2 s 387982 0 388038 800 6 la_data_out[80]
port 378 nsew signal output
rlabel metal2 s 391294 0 391350 800 6 la_data_out[81]
port 379 nsew signal output
rlabel metal2 s 394606 0 394662 800 6 la_data_out[82]
port 380 nsew signal output
rlabel metal2 s 397918 0 397974 800 6 la_data_out[83]
port 381 nsew signal output
rlabel metal2 s 401230 0 401286 800 6 la_data_out[84]
port 382 nsew signal output
rlabel metal2 s 404542 0 404598 800 6 la_data_out[85]
port 383 nsew signal output
rlabel metal2 s 407854 0 407910 800 6 la_data_out[86]
port 384 nsew signal output
rlabel metal2 s 411166 0 411222 800 6 la_data_out[87]
port 385 nsew signal output
rlabel metal2 s 414478 0 414534 800 6 la_data_out[88]
port 386 nsew signal output
rlabel metal2 s 417790 0 417846 800 6 la_data_out[89]
port 387 nsew signal output
rlabel metal2 s 149518 0 149574 800 6 la_data_out[8]
port 388 nsew signal output
rlabel metal2 s 421102 0 421158 800 6 la_data_out[90]
port 389 nsew signal output
rlabel metal2 s 424414 0 424470 800 6 la_data_out[91]
port 390 nsew signal output
rlabel metal2 s 427726 0 427782 800 6 la_data_out[92]
port 391 nsew signal output
rlabel metal2 s 431038 0 431094 800 6 la_data_out[93]
port 392 nsew signal output
rlabel metal2 s 434350 0 434406 800 6 la_data_out[94]
port 393 nsew signal output
rlabel metal2 s 437662 0 437718 800 6 la_data_out[95]
port 394 nsew signal output
rlabel metal2 s 440974 0 441030 800 6 la_data_out[96]
port 395 nsew signal output
rlabel metal2 s 444286 0 444342 800 6 la_data_out[97]
port 396 nsew signal output
rlabel metal2 s 447598 0 447654 800 6 la_data_out[98]
port 397 nsew signal output
rlabel metal2 s 450910 0 450966 800 6 la_data_out[99]
port 398 nsew signal output
rlabel metal2 s 152830 0 152886 800 6 la_data_out[9]
port 399 nsew signal output
rlabel metal2 s 124126 0 124182 800 6 la_oenb[0]
port 400 nsew signal input
rlabel metal2 s 455326 0 455382 800 6 la_oenb[100]
port 401 nsew signal input
rlabel metal2 s 458638 0 458694 800 6 la_oenb[101]
port 402 nsew signal input
rlabel metal2 s 461950 0 462006 800 6 la_oenb[102]
port 403 nsew signal input
rlabel metal2 s 465262 0 465318 800 6 la_oenb[103]
port 404 nsew signal input
rlabel metal2 s 468574 0 468630 800 6 la_oenb[104]
port 405 nsew signal input
rlabel metal2 s 471886 0 471942 800 6 la_oenb[105]
port 406 nsew signal input
rlabel metal2 s 475198 0 475254 800 6 la_oenb[106]
port 407 nsew signal input
rlabel metal2 s 478510 0 478566 800 6 la_oenb[107]
port 408 nsew signal input
rlabel metal2 s 481822 0 481878 800 6 la_oenb[108]
port 409 nsew signal input
rlabel metal2 s 485134 0 485190 800 6 la_oenb[109]
port 410 nsew signal input
rlabel metal2 s 157246 0 157302 800 6 la_oenb[10]
port 411 nsew signal input
rlabel metal2 s 488446 0 488502 800 6 la_oenb[110]
port 412 nsew signal input
rlabel metal2 s 491758 0 491814 800 6 la_oenb[111]
port 413 nsew signal input
rlabel metal2 s 495070 0 495126 800 6 la_oenb[112]
port 414 nsew signal input
rlabel metal2 s 498382 0 498438 800 6 la_oenb[113]
port 415 nsew signal input
rlabel metal2 s 501694 0 501750 800 6 la_oenb[114]
port 416 nsew signal input
rlabel metal2 s 505006 0 505062 800 6 la_oenb[115]
port 417 nsew signal input
rlabel metal2 s 508318 0 508374 800 6 la_oenb[116]
port 418 nsew signal input
rlabel metal2 s 511630 0 511686 800 6 la_oenb[117]
port 419 nsew signal input
rlabel metal2 s 514942 0 514998 800 6 la_oenb[118]
port 420 nsew signal input
rlabel metal2 s 518254 0 518310 800 6 la_oenb[119]
port 421 nsew signal input
rlabel metal2 s 160558 0 160614 800 6 la_oenb[11]
port 422 nsew signal input
rlabel metal2 s 521566 0 521622 800 6 la_oenb[120]
port 423 nsew signal input
rlabel metal2 s 524878 0 524934 800 6 la_oenb[121]
port 424 nsew signal input
rlabel metal2 s 528190 0 528246 800 6 la_oenb[122]
port 425 nsew signal input
rlabel metal2 s 531502 0 531558 800 6 la_oenb[123]
port 426 nsew signal input
rlabel metal2 s 534814 0 534870 800 6 la_oenb[124]
port 427 nsew signal input
rlabel metal2 s 538126 0 538182 800 6 la_oenb[125]
port 428 nsew signal input
rlabel metal2 s 541438 0 541494 800 6 la_oenb[126]
port 429 nsew signal input
rlabel metal2 s 544750 0 544806 800 6 la_oenb[127]
port 430 nsew signal input
rlabel metal2 s 163870 0 163926 800 6 la_oenb[12]
port 431 nsew signal input
rlabel metal2 s 167182 0 167238 800 6 la_oenb[13]
port 432 nsew signal input
rlabel metal2 s 170494 0 170550 800 6 la_oenb[14]
port 433 nsew signal input
rlabel metal2 s 173806 0 173862 800 6 la_oenb[15]
port 434 nsew signal input
rlabel metal2 s 177118 0 177174 800 6 la_oenb[16]
port 435 nsew signal input
rlabel metal2 s 180430 0 180486 800 6 la_oenb[17]
port 436 nsew signal input
rlabel metal2 s 183742 0 183798 800 6 la_oenb[18]
port 437 nsew signal input
rlabel metal2 s 187054 0 187110 800 6 la_oenb[19]
port 438 nsew signal input
rlabel metal2 s 127438 0 127494 800 6 la_oenb[1]
port 439 nsew signal input
rlabel metal2 s 190366 0 190422 800 6 la_oenb[20]
port 440 nsew signal input
rlabel metal2 s 193678 0 193734 800 6 la_oenb[21]
port 441 nsew signal input
rlabel metal2 s 196990 0 197046 800 6 la_oenb[22]
port 442 nsew signal input
rlabel metal2 s 200302 0 200358 800 6 la_oenb[23]
port 443 nsew signal input
rlabel metal2 s 203614 0 203670 800 6 la_oenb[24]
port 444 nsew signal input
rlabel metal2 s 206926 0 206982 800 6 la_oenb[25]
port 445 nsew signal input
rlabel metal2 s 210238 0 210294 800 6 la_oenb[26]
port 446 nsew signal input
rlabel metal2 s 213550 0 213606 800 6 la_oenb[27]
port 447 nsew signal input
rlabel metal2 s 216862 0 216918 800 6 la_oenb[28]
port 448 nsew signal input
rlabel metal2 s 220174 0 220230 800 6 la_oenb[29]
port 449 nsew signal input
rlabel metal2 s 130750 0 130806 800 6 la_oenb[2]
port 450 nsew signal input
rlabel metal2 s 223486 0 223542 800 6 la_oenb[30]
port 451 nsew signal input
rlabel metal2 s 226798 0 226854 800 6 la_oenb[31]
port 452 nsew signal input
rlabel metal2 s 230110 0 230166 800 6 la_oenb[32]
port 453 nsew signal input
rlabel metal2 s 233422 0 233478 800 6 la_oenb[33]
port 454 nsew signal input
rlabel metal2 s 236734 0 236790 800 6 la_oenb[34]
port 455 nsew signal input
rlabel metal2 s 240046 0 240102 800 6 la_oenb[35]
port 456 nsew signal input
rlabel metal2 s 243358 0 243414 800 6 la_oenb[36]
port 457 nsew signal input
rlabel metal2 s 246670 0 246726 800 6 la_oenb[37]
port 458 nsew signal input
rlabel metal2 s 249982 0 250038 800 6 la_oenb[38]
port 459 nsew signal input
rlabel metal2 s 253294 0 253350 800 6 la_oenb[39]
port 460 nsew signal input
rlabel metal2 s 134062 0 134118 800 6 la_oenb[3]
port 461 nsew signal input
rlabel metal2 s 256606 0 256662 800 6 la_oenb[40]
port 462 nsew signal input
rlabel metal2 s 259918 0 259974 800 6 la_oenb[41]
port 463 nsew signal input
rlabel metal2 s 263230 0 263286 800 6 la_oenb[42]
port 464 nsew signal input
rlabel metal2 s 266542 0 266598 800 6 la_oenb[43]
port 465 nsew signal input
rlabel metal2 s 269854 0 269910 800 6 la_oenb[44]
port 466 nsew signal input
rlabel metal2 s 273166 0 273222 800 6 la_oenb[45]
port 467 nsew signal input
rlabel metal2 s 276478 0 276534 800 6 la_oenb[46]
port 468 nsew signal input
rlabel metal2 s 279790 0 279846 800 6 la_oenb[47]
port 469 nsew signal input
rlabel metal2 s 283102 0 283158 800 6 la_oenb[48]
port 470 nsew signal input
rlabel metal2 s 286414 0 286470 800 6 la_oenb[49]
port 471 nsew signal input
rlabel metal2 s 137374 0 137430 800 6 la_oenb[4]
port 472 nsew signal input
rlabel metal2 s 289726 0 289782 800 6 la_oenb[50]
port 473 nsew signal input
rlabel metal2 s 293038 0 293094 800 6 la_oenb[51]
port 474 nsew signal input
rlabel metal2 s 296350 0 296406 800 6 la_oenb[52]
port 475 nsew signal input
rlabel metal2 s 299662 0 299718 800 6 la_oenb[53]
port 476 nsew signal input
rlabel metal2 s 302974 0 303030 800 6 la_oenb[54]
port 477 nsew signal input
rlabel metal2 s 306286 0 306342 800 6 la_oenb[55]
port 478 nsew signal input
rlabel metal2 s 309598 0 309654 800 6 la_oenb[56]
port 479 nsew signal input
rlabel metal2 s 312910 0 312966 800 6 la_oenb[57]
port 480 nsew signal input
rlabel metal2 s 316222 0 316278 800 6 la_oenb[58]
port 481 nsew signal input
rlabel metal2 s 319534 0 319590 800 6 la_oenb[59]
port 482 nsew signal input
rlabel metal2 s 140686 0 140742 800 6 la_oenb[5]
port 483 nsew signal input
rlabel metal2 s 322846 0 322902 800 6 la_oenb[60]
port 484 nsew signal input
rlabel metal2 s 326158 0 326214 800 6 la_oenb[61]
port 485 nsew signal input
rlabel metal2 s 329470 0 329526 800 6 la_oenb[62]
port 486 nsew signal input
rlabel metal2 s 332782 0 332838 800 6 la_oenb[63]
port 487 nsew signal input
rlabel metal2 s 336094 0 336150 800 6 la_oenb[64]
port 488 nsew signal input
rlabel metal2 s 339406 0 339462 800 6 la_oenb[65]
port 489 nsew signal input
rlabel metal2 s 342718 0 342774 800 6 la_oenb[66]
port 490 nsew signal input
rlabel metal2 s 346030 0 346086 800 6 la_oenb[67]
port 491 nsew signal input
rlabel metal2 s 349342 0 349398 800 6 la_oenb[68]
port 492 nsew signal input
rlabel metal2 s 352654 0 352710 800 6 la_oenb[69]
port 493 nsew signal input
rlabel metal2 s 143998 0 144054 800 6 la_oenb[6]
port 494 nsew signal input
rlabel metal2 s 355966 0 356022 800 6 la_oenb[70]
port 495 nsew signal input
rlabel metal2 s 359278 0 359334 800 6 la_oenb[71]
port 496 nsew signal input
rlabel metal2 s 362590 0 362646 800 6 la_oenb[72]
port 497 nsew signal input
rlabel metal2 s 365902 0 365958 800 6 la_oenb[73]
port 498 nsew signal input
rlabel metal2 s 369214 0 369270 800 6 la_oenb[74]
port 499 nsew signal input
rlabel metal2 s 372526 0 372582 800 6 la_oenb[75]
port 500 nsew signal input
rlabel metal2 s 375838 0 375894 800 6 la_oenb[76]
port 501 nsew signal input
rlabel metal2 s 379150 0 379206 800 6 la_oenb[77]
port 502 nsew signal input
rlabel metal2 s 382462 0 382518 800 6 la_oenb[78]
port 503 nsew signal input
rlabel metal2 s 385774 0 385830 800 6 la_oenb[79]
port 504 nsew signal input
rlabel metal2 s 147310 0 147366 800 6 la_oenb[7]
port 505 nsew signal input
rlabel metal2 s 389086 0 389142 800 6 la_oenb[80]
port 506 nsew signal input
rlabel metal2 s 392398 0 392454 800 6 la_oenb[81]
port 507 nsew signal input
rlabel metal2 s 395710 0 395766 800 6 la_oenb[82]
port 508 nsew signal input
rlabel metal2 s 399022 0 399078 800 6 la_oenb[83]
port 509 nsew signal input
rlabel metal2 s 402334 0 402390 800 6 la_oenb[84]
port 510 nsew signal input
rlabel metal2 s 405646 0 405702 800 6 la_oenb[85]
port 511 nsew signal input
rlabel metal2 s 408958 0 409014 800 6 la_oenb[86]
port 512 nsew signal input
rlabel metal2 s 412270 0 412326 800 6 la_oenb[87]
port 513 nsew signal input
rlabel metal2 s 415582 0 415638 800 6 la_oenb[88]
port 514 nsew signal input
rlabel metal2 s 418894 0 418950 800 6 la_oenb[89]
port 515 nsew signal input
rlabel metal2 s 150622 0 150678 800 6 la_oenb[8]
port 516 nsew signal input
rlabel metal2 s 422206 0 422262 800 6 la_oenb[90]
port 517 nsew signal input
rlabel metal2 s 425518 0 425574 800 6 la_oenb[91]
port 518 nsew signal input
rlabel metal2 s 428830 0 428886 800 6 la_oenb[92]
port 519 nsew signal input
rlabel metal2 s 432142 0 432198 800 6 la_oenb[93]
port 520 nsew signal input
rlabel metal2 s 435454 0 435510 800 6 la_oenb[94]
port 521 nsew signal input
rlabel metal2 s 438766 0 438822 800 6 la_oenb[95]
port 522 nsew signal input
rlabel metal2 s 442078 0 442134 800 6 la_oenb[96]
port 523 nsew signal input
rlabel metal2 s 445390 0 445446 800 6 la_oenb[97]
port 524 nsew signal input
rlabel metal2 s 448702 0 448758 800 6 la_oenb[98]
port 525 nsew signal input
rlabel metal2 s 452014 0 452070 800 6 la_oenb[99]
port 526 nsew signal input
rlabel metal2 s 153934 0 153990 800 6 la_oenb[9]
port 527 nsew signal input
rlabel metal2 s 545854 0 545910 800 6 user_clock2
port 528 nsew signal input
rlabel metal2 s 546958 0 547014 800 6 user_irq[0]
port 529 nsew signal output
rlabel metal2 s 548062 0 548118 800 6 user_irq[1]
port 530 nsew signal output
rlabel metal2 s 549166 0 549222 800 6 user_irq[2]
port 531 nsew signal output
rlabel metal4 s 4208 2128 4528 664272 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 664272 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 664272 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 664272 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 664272 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 664272 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 188528 2128 188848 664272 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 219248 2128 219568 664272 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 249968 2128 250288 664272 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 280688 2128 281008 664272 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 311408 2128 311728 664272 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 342128 2128 342448 664272 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 372848 2128 373168 664272 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 403568 2128 403888 664272 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 434288 2128 434608 664272 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 465008 2128 465328 664272 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 495728 2128 496048 664272 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 526448 2128 526768 664272 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 664272 6 vssd1
port 533 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 664272 6 vssd1
port 533 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 664272 6 vssd1
port 533 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 664272 6 vssd1
port 533 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 664272 6 vssd1
port 533 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 664272 6 vssd1
port 533 nsew ground bidirectional
rlabel metal4 s 203888 2128 204208 664272 6 vssd1
port 533 nsew ground bidirectional
rlabel metal4 s 234608 2128 234928 664272 6 vssd1
port 533 nsew ground bidirectional
rlabel metal4 s 265328 2128 265648 664272 6 vssd1
port 533 nsew ground bidirectional
rlabel metal4 s 296048 2128 296368 664272 6 vssd1
port 533 nsew ground bidirectional
rlabel metal4 s 326768 2128 327088 664272 6 vssd1
port 533 nsew ground bidirectional
rlabel metal4 s 357488 2128 357808 664272 6 vssd1
port 533 nsew ground bidirectional
rlabel metal4 s 388208 2128 388528 664272 6 vssd1
port 533 nsew ground bidirectional
rlabel metal4 s 418928 2128 419248 664272 6 vssd1
port 533 nsew ground bidirectional
rlabel metal4 s 449648 2128 449968 664272 6 vssd1
port 533 nsew ground bidirectional
rlabel metal4 s 480368 2128 480688 664272 6 vssd1
port 533 nsew ground bidirectional
rlabel metal4 s 511088 2128 511408 664272 6 vssd1
port 533 nsew ground bidirectional
rlabel metal4 s 541808 2128 542128 664272 6 vssd1
port 533 nsew ground bidirectional
rlabel metal2 s 4894 0 4950 800 6 wb_clk_i
port 534 nsew signal input
rlabel metal2 s 5998 0 6054 800 6 wb_rst_i
port 535 nsew signal input
rlabel metal2 s 7102 0 7158 800 6 wbs_ack_o
port 536 nsew signal output
rlabel metal2 s 11518 0 11574 800 6 wbs_adr_i[0]
port 537 nsew signal input
rlabel metal2 s 49054 0 49110 800 6 wbs_adr_i[10]
port 538 nsew signal input
rlabel metal2 s 52366 0 52422 800 6 wbs_adr_i[11]
port 539 nsew signal input
rlabel metal2 s 55678 0 55734 800 6 wbs_adr_i[12]
port 540 nsew signal input
rlabel metal2 s 58990 0 59046 800 6 wbs_adr_i[13]
port 541 nsew signal input
rlabel metal2 s 62302 0 62358 800 6 wbs_adr_i[14]
port 542 nsew signal input
rlabel metal2 s 65614 0 65670 800 6 wbs_adr_i[15]
port 543 nsew signal input
rlabel metal2 s 68926 0 68982 800 6 wbs_adr_i[16]
port 544 nsew signal input
rlabel metal2 s 72238 0 72294 800 6 wbs_adr_i[17]
port 545 nsew signal input
rlabel metal2 s 75550 0 75606 800 6 wbs_adr_i[18]
port 546 nsew signal input
rlabel metal2 s 78862 0 78918 800 6 wbs_adr_i[19]
port 547 nsew signal input
rlabel metal2 s 15934 0 15990 800 6 wbs_adr_i[1]
port 548 nsew signal input
rlabel metal2 s 82174 0 82230 800 6 wbs_adr_i[20]
port 549 nsew signal input
rlabel metal2 s 85486 0 85542 800 6 wbs_adr_i[21]
port 550 nsew signal input
rlabel metal2 s 88798 0 88854 800 6 wbs_adr_i[22]
port 551 nsew signal input
rlabel metal2 s 92110 0 92166 800 6 wbs_adr_i[23]
port 552 nsew signal input
rlabel metal2 s 95422 0 95478 800 6 wbs_adr_i[24]
port 553 nsew signal input
rlabel metal2 s 98734 0 98790 800 6 wbs_adr_i[25]
port 554 nsew signal input
rlabel metal2 s 102046 0 102102 800 6 wbs_adr_i[26]
port 555 nsew signal input
rlabel metal2 s 105358 0 105414 800 6 wbs_adr_i[27]
port 556 nsew signal input
rlabel metal2 s 108670 0 108726 800 6 wbs_adr_i[28]
port 557 nsew signal input
rlabel metal2 s 111982 0 112038 800 6 wbs_adr_i[29]
port 558 nsew signal input
rlabel metal2 s 20350 0 20406 800 6 wbs_adr_i[2]
port 559 nsew signal input
rlabel metal2 s 115294 0 115350 800 6 wbs_adr_i[30]
port 560 nsew signal input
rlabel metal2 s 118606 0 118662 800 6 wbs_adr_i[31]
port 561 nsew signal input
rlabel metal2 s 24766 0 24822 800 6 wbs_adr_i[3]
port 562 nsew signal input
rlabel metal2 s 29182 0 29238 800 6 wbs_adr_i[4]
port 563 nsew signal input
rlabel metal2 s 32494 0 32550 800 6 wbs_adr_i[5]
port 564 nsew signal input
rlabel metal2 s 35806 0 35862 800 6 wbs_adr_i[6]
port 565 nsew signal input
rlabel metal2 s 39118 0 39174 800 6 wbs_adr_i[7]
port 566 nsew signal input
rlabel metal2 s 42430 0 42486 800 6 wbs_adr_i[8]
port 567 nsew signal input
rlabel metal2 s 45742 0 45798 800 6 wbs_adr_i[9]
port 568 nsew signal input
rlabel metal2 s 8206 0 8262 800 6 wbs_cyc_i
port 569 nsew signal input
rlabel metal2 s 12622 0 12678 800 6 wbs_dat_i[0]
port 570 nsew signal input
rlabel metal2 s 50158 0 50214 800 6 wbs_dat_i[10]
port 571 nsew signal input
rlabel metal2 s 53470 0 53526 800 6 wbs_dat_i[11]
port 572 nsew signal input
rlabel metal2 s 56782 0 56838 800 6 wbs_dat_i[12]
port 573 nsew signal input
rlabel metal2 s 60094 0 60150 800 6 wbs_dat_i[13]
port 574 nsew signal input
rlabel metal2 s 63406 0 63462 800 6 wbs_dat_i[14]
port 575 nsew signal input
rlabel metal2 s 66718 0 66774 800 6 wbs_dat_i[15]
port 576 nsew signal input
rlabel metal2 s 70030 0 70086 800 6 wbs_dat_i[16]
port 577 nsew signal input
rlabel metal2 s 73342 0 73398 800 6 wbs_dat_i[17]
port 578 nsew signal input
rlabel metal2 s 76654 0 76710 800 6 wbs_dat_i[18]
port 579 nsew signal input
rlabel metal2 s 79966 0 80022 800 6 wbs_dat_i[19]
port 580 nsew signal input
rlabel metal2 s 17038 0 17094 800 6 wbs_dat_i[1]
port 581 nsew signal input
rlabel metal2 s 83278 0 83334 800 6 wbs_dat_i[20]
port 582 nsew signal input
rlabel metal2 s 86590 0 86646 800 6 wbs_dat_i[21]
port 583 nsew signal input
rlabel metal2 s 89902 0 89958 800 6 wbs_dat_i[22]
port 584 nsew signal input
rlabel metal2 s 93214 0 93270 800 6 wbs_dat_i[23]
port 585 nsew signal input
rlabel metal2 s 96526 0 96582 800 6 wbs_dat_i[24]
port 586 nsew signal input
rlabel metal2 s 99838 0 99894 800 6 wbs_dat_i[25]
port 587 nsew signal input
rlabel metal2 s 103150 0 103206 800 6 wbs_dat_i[26]
port 588 nsew signal input
rlabel metal2 s 106462 0 106518 800 6 wbs_dat_i[27]
port 589 nsew signal input
rlabel metal2 s 109774 0 109830 800 6 wbs_dat_i[28]
port 590 nsew signal input
rlabel metal2 s 113086 0 113142 800 6 wbs_dat_i[29]
port 591 nsew signal input
rlabel metal2 s 21454 0 21510 800 6 wbs_dat_i[2]
port 592 nsew signal input
rlabel metal2 s 116398 0 116454 800 6 wbs_dat_i[30]
port 593 nsew signal input
rlabel metal2 s 119710 0 119766 800 6 wbs_dat_i[31]
port 594 nsew signal input
rlabel metal2 s 25870 0 25926 800 6 wbs_dat_i[3]
port 595 nsew signal input
rlabel metal2 s 30286 0 30342 800 6 wbs_dat_i[4]
port 596 nsew signal input
rlabel metal2 s 33598 0 33654 800 6 wbs_dat_i[5]
port 597 nsew signal input
rlabel metal2 s 36910 0 36966 800 6 wbs_dat_i[6]
port 598 nsew signal input
rlabel metal2 s 40222 0 40278 800 6 wbs_dat_i[7]
port 599 nsew signal input
rlabel metal2 s 43534 0 43590 800 6 wbs_dat_i[8]
port 600 nsew signal input
rlabel metal2 s 46846 0 46902 800 6 wbs_dat_i[9]
port 601 nsew signal input
rlabel metal2 s 13726 0 13782 800 6 wbs_dat_o[0]
port 602 nsew signal output
rlabel metal2 s 51262 0 51318 800 6 wbs_dat_o[10]
port 603 nsew signal output
rlabel metal2 s 54574 0 54630 800 6 wbs_dat_o[11]
port 604 nsew signal output
rlabel metal2 s 57886 0 57942 800 6 wbs_dat_o[12]
port 605 nsew signal output
rlabel metal2 s 61198 0 61254 800 6 wbs_dat_o[13]
port 606 nsew signal output
rlabel metal2 s 64510 0 64566 800 6 wbs_dat_o[14]
port 607 nsew signal output
rlabel metal2 s 67822 0 67878 800 6 wbs_dat_o[15]
port 608 nsew signal output
rlabel metal2 s 71134 0 71190 800 6 wbs_dat_o[16]
port 609 nsew signal output
rlabel metal2 s 74446 0 74502 800 6 wbs_dat_o[17]
port 610 nsew signal output
rlabel metal2 s 77758 0 77814 800 6 wbs_dat_o[18]
port 611 nsew signal output
rlabel metal2 s 81070 0 81126 800 6 wbs_dat_o[19]
port 612 nsew signal output
rlabel metal2 s 18142 0 18198 800 6 wbs_dat_o[1]
port 613 nsew signal output
rlabel metal2 s 84382 0 84438 800 6 wbs_dat_o[20]
port 614 nsew signal output
rlabel metal2 s 87694 0 87750 800 6 wbs_dat_o[21]
port 615 nsew signal output
rlabel metal2 s 91006 0 91062 800 6 wbs_dat_o[22]
port 616 nsew signal output
rlabel metal2 s 94318 0 94374 800 6 wbs_dat_o[23]
port 617 nsew signal output
rlabel metal2 s 97630 0 97686 800 6 wbs_dat_o[24]
port 618 nsew signal output
rlabel metal2 s 100942 0 100998 800 6 wbs_dat_o[25]
port 619 nsew signal output
rlabel metal2 s 104254 0 104310 800 6 wbs_dat_o[26]
port 620 nsew signal output
rlabel metal2 s 107566 0 107622 800 6 wbs_dat_o[27]
port 621 nsew signal output
rlabel metal2 s 110878 0 110934 800 6 wbs_dat_o[28]
port 622 nsew signal output
rlabel metal2 s 114190 0 114246 800 6 wbs_dat_o[29]
port 623 nsew signal output
rlabel metal2 s 22558 0 22614 800 6 wbs_dat_o[2]
port 624 nsew signal output
rlabel metal2 s 117502 0 117558 800 6 wbs_dat_o[30]
port 625 nsew signal output
rlabel metal2 s 120814 0 120870 800 6 wbs_dat_o[31]
port 626 nsew signal output
rlabel metal2 s 26974 0 27030 800 6 wbs_dat_o[3]
port 627 nsew signal output
rlabel metal2 s 31390 0 31446 800 6 wbs_dat_o[4]
port 628 nsew signal output
rlabel metal2 s 34702 0 34758 800 6 wbs_dat_o[5]
port 629 nsew signal output
rlabel metal2 s 38014 0 38070 800 6 wbs_dat_o[6]
port 630 nsew signal output
rlabel metal2 s 41326 0 41382 800 6 wbs_dat_o[7]
port 631 nsew signal output
rlabel metal2 s 44638 0 44694 800 6 wbs_dat_o[8]
port 632 nsew signal output
rlabel metal2 s 47950 0 48006 800 6 wbs_dat_o[9]
port 633 nsew signal output
rlabel metal2 s 14830 0 14886 800 6 wbs_sel_i[0]
port 634 nsew signal input
rlabel metal2 s 19246 0 19302 800 6 wbs_sel_i[1]
port 635 nsew signal input
rlabel metal2 s 23662 0 23718 800 6 wbs_sel_i[2]
port 636 nsew signal input
rlabel metal2 s 28078 0 28134 800 6 wbs_sel_i[3]
port 637 nsew signal input
rlabel metal2 s 9310 0 9366 800 6 wbs_stb_i
port 638 nsew signal input
rlabel metal2 s 10414 0 10470 800 6 wbs_we_i
port 639 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 554204 666748
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 800896442
string GDS_FILE /mnt/r/work/Rift2Go_2320_Sky130_MPW8/openlane/user_proj_example/runs/22_11_23_20_50/results/signoff/rift2Wrap.magic.gds
string GDS_START 2039606
<< end >>

